
#******
# Preview export LEF
#
#	 Preview sub-version 5.10.41.500.0.10
#
# TECH LIB NAME: ts018_prim
# TECH FILE NAME: techfile.cds
#******

VERSION 5.4 ;

NAMESCASESENSITIVE ON ;

DIVIDERCHAR "/" ;
BUSBITCHARS "[]" ;

UNITS
    DATABASE MICRONS 1000  ;
END UNITS

 MANUFACTURINGGRID    0.005000 ;

SITE IOSite_c
    SYMMETRY X Y  R90   ;
    CLASS PAD  ;
    SIZE 0.010 BY 250.000 ;
END IOSite_c

SITE CO_MSTR_c
        CLASS PAD ;
        SIZE  250.000 BY 250.000 ;
END CO_MSTR_c

MACRO pvdi
    CLASS PAD ;
    FOREIGN pvdi 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 65.000 BY 250.000 ;
    SYMMETRY X Y R90 ;
    SITE IOSite_c ;
    PIN VDDO
        DIRECTION INOUT ;
        USE power ;
        PORT
        LAYER M3 ;
        RECT  64.200 192.330 65.000 200.640 ;
        RECT  0.000 201.660 65.000 221.520 ;
        RECT  0.000 222.720 65.000 246.820 ;
        RECT  0.000 192.330 0.800 200.640 ;
        LAYER M2 ;
        RECT  0.000 186.470 65.000 195.650 ;
        LAYER TOP_M ;
        RECT  62.900 195.170 65.000 200.640 ;
        RECT  62.900 201.660 65.000 221.520 ;
        RECT  62.900 222.720 65.000 246.820 ;
        RECT  0.000 195.170 2.100 200.640 ;
        RECT  0.000 201.660 2.100 221.520 ;
        RECT  0.000 222.720 2.100 246.820 ;
        END
    END VDDO
    PIN VDD
        DIRECTION OUTPUT ;
        USE power ;
        PORT
	CLASS CORE ;
        LAYER M3 ;
        RECT  64.200 163.510 65.000 190.890 ;
        RECT  15.560 247.440 49.380 250.000 ;
        RECT  0.000 163.510 0.800 190.890 ;
        LAYER M2 ;
        RECT  0.000 172.080 65.000 183.060 ;
        RECT  2.000 61.000 63.000 90.230 ;
        RECT  15.560 246.600 49.380 250.000 ;
        LAYER TOP_M ;
        RECT  62.900 163.500 65.000 194.560 ;
        RECT  15.560 247.440 49.380 250.000 ;
        RECT  0.000 163.500 2.100 194.560 ;
        END
    END VDD
    PIN VSSO
        DIRECTION INOUT ;
        USE ground ;
        PORT
        LAYER M3 ;
        RECT  0.000 92.060 65.000 123.250 ;
        RECT  64.200 149.940 65.000 162.610 ;
        RECT  0.000 149.940 0.800 162.610 ;
        LAYER M2 ;
        RECT  0.000 147.040 65.000 154.520 ;
        LAYER TOP_M ;
        RECT  62.900 92.060 65.000 123.250 ;
        RECT  62.900 155.410 65.000 162.610 ;
        RECT  0.000 92.060 2.100 123.250 ;
        RECT  0.000 155.410 2.100 162.610 ;
        END
    END VSSO
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        PORT
        LAYER M3 ;
        RECT  64.200 130.690 65.000 148.880 ;
        RECT  0.000 130.690 0.800 148.880 ;
        LAYER M2 ;
        RECT  0.000 136.310 65.000 146.340 ;
        LAYER TOP_M ;
        RECT  62.900 123.850 65.000 154.560 ;
        RECT  0.000 123.850 2.100 154.560 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  2.000 0.000 63.000 250.000 ;
        RECT  0.000 88.990 65.000 130.360 ;
        RECT  0.000 136.510 65.000 157.550 ;
        RECT  0.500 136.510 64.500 163.550 ;
        RECT  0.600 0.600 64.400 250.000 ;
        RECT  0.000 198.470 65.000 250.000 ;
        LAYER M2 ;
        RECT  0.600 196.440 64.400 245.810 ;
        RECT  12.630 196.340 14.950 246.720 ;
        RECT  50.060 196.440 64.400 246.720 ;
        RECT  0.600 196.440 14.770 249.400 ;
        RECT  50.170 196.440 64.400 249.400 ;
        RECT  0.600 183.850 64.400 185.680 ;
        RECT  0.600 155.310 64.400 171.290 ;
        RECT  2.000 0.000 63.000 60.210 ;
        RECT  0.600 0.600 64.400 60.210 ;
        RECT  0.600 0.600 1.210 135.520 ;
        RECT  0.600 91.020 64.400 135.520 ;
        RECT  4.080 91.020 60.940 135.690 ;
        LAYER M3 ;
        RECT  0.600 247.660 14.720 249.400 ;
        RECT  50.220 247.660 64.400 249.400 ;
        RECT  0.600 0.600 64.400 60.480 ;
        RECT  2.000 0.000 63.000 88.700 ;
        RECT  0.600 0.600 1.480 91.220 ;
        RECT  0.600 90.750 64.400 91.220 ;
        RECT  0.600 124.090 64.650 128.560 ;
        RECT  0.600 124.090 64.400 129.850 ;
        RECT  1.400 124.090 63.595 135.790 ;
        RECT  3.070 124.090 58.100 200.820 ;
        RECT  62.470 124.090 63.595 154.120 ;
        RECT  1.400 124.090 2.470 154.470 ;
        RECT  1.640 155.040 63.360 171.560 ;
        RECT  1.640 183.580 63.360 185.950 ;
        RECT  3.070 144.980 61.290 200.820 ;
        RECT  1.640 196.170 63.360 200.820 ;
        RECT  58.010 144.980 59.020 201.060 ;
        RECT  60.060 144.980 61.290 201.060 ;
        LAYER TOP_M ;
        RECT  2.970 247.550 14.690 249.400 ;
        RECT  0.600 247.690 14.690 249.400 ;
        RECT  2.970 222.720 62.030 246.820 ;
        RECT  2.970 201.660 62.030 221.520 ;
        RECT  2.970 123.850 62.030 200.930 ;
        RECT  2.970 92.060 62.030 123.250 ;
        RECT  50.250 247.550 62.030 249.400 ;
        RECT  50.250 247.690 64.400 249.400 ;
        RECT  2.000 0.000 63.000 91.190 ;
        RECT  0.600 0.600 64.400 91.190 ;
        RECT  2.970 0.000 62.030 91.330 ;
    END
END pvdi

MACRO pvdc
    CLASS PAD ;
    FOREIGN pvdc 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 65.000 BY 250.000 ;
    SYMMETRY X Y R90 ;
    SITE IOSite_c ;
    PIN VDDO
        DIRECTION INOUT ;
        USE power ;
        PORT
        LAYER M3 ;
        RECT  64.200 192.330 65.000 200.640 ;
        RECT  0.000 201.660 65.000 221.520 ;
        RECT  0.000 222.720 65.000 246.820 ;
        RECT  0.000 192.330 0.800 200.640 ;
        LAYER M2 ;
        RECT  0.000 186.470 65.000 195.650 ;
        LAYER TOP_M ;
        RECT  62.900 195.170 65.000 200.640 ;
        RECT  62.900 201.660 65.000 221.520 ;
        RECT  62.900 222.720 65.000 246.820 ;
        RECT  0.000 195.170 2.100 200.640 ;
        RECT  0.000 201.660 2.100 221.520 ;
        RECT  0.000 222.720 2.100 246.820 ;
        END
    END VDDO
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        PORT
        LAYER M3 ;
        RECT  64.200 163.510 65.000 190.890 ;
        RECT  0.000 163.510 0.800 190.890 ;
        LAYER M2 ;
        RECT  0.000 172.080 65.000 183.060 ;
        LAYER TOP_M ;
        RECT  62.900 163.500 65.000 194.560 ;
        RECT  0.000 163.500 2.100 194.560 ;
        END
    END VDD
    PIN VSSO
        DIRECTION INOUT ;
        USE ground ;
        PORT
        LAYER M3 ;
        RECT  0.000 92.060 65.000 123.250 ;
        RECT  64.200 149.940 65.000 162.610 ;
        RECT  0.000 149.940 0.800 162.610 ;
        LAYER M2 ;
        RECT  0.000 147.040 65.000 154.520 ;
        LAYER TOP_M ;
        RECT  62.900 92.060 65.000 123.250 ;
        RECT  62.900 155.410 65.000 162.610 ;
        RECT  0.000 92.060 2.100 123.250 ;
        RECT  0.000 155.410 2.100 162.610 ;
        END
    END VSSO
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        PORT
        LAYER M3 ;
        RECT  64.200 130.690 65.000 148.880 ;
        RECT  0.000 130.690 0.800 148.880 ;
        LAYER M2 ;
        RECT  0.000 136.310 65.000 146.340 ;
        LAYER TOP_M ;
        RECT  62.900 123.850 65.000 154.560 ;
        RECT  0.000 123.850 2.100 154.560 ;
        END
    END VSS
    PIN VDDC
        DIRECTION OUTPUT ;
        USE power ;
        PORT
	CLASS CORE ;
        LAYER M3 ;
        RECT  15.560 247.710 49.380 250.000 ;
        LAYER M2 ;
        RECT  2.000 61.000 63.000 90.230 ;
        RECT  15.560 246.120 49.380 250.000 ;
        LAYER TOP_M ;
        RECT  15.560 247.420 49.380 250.000 ;
        END
    END VDDC
    OBS
        LAYER M1 ;
        RECT  2.000 0.000 63.000 250.000 ;
        RECT  0.000 88.990 65.000 130.360 ;
        RECT  0.000 136.510 65.000 157.550 ;
        RECT  0.500 136.510 64.500 163.550 ;
        RECT  0.600 0.600 64.400 250.000 ;
        RECT  0.000 198.470 65.000 250.000 ;
        LAYER M2 ;
        RECT  0.600 196.440 64.400 245.330 ;
        RECT  12.640 196.370 14.950 246.720 ;
        RECT  50.060 196.440 64.400 246.720 ;
        RECT  0.600 196.440 14.770 249.400 ;
        RECT  50.170 196.440 64.400 249.400 ;
        RECT  0.600 183.850 64.400 185.680 ;
        RECT  0.600 155.310 64.400 171.290 ;
        RECT  2.000 0.000 63.000 60.210 ;
        RECT  0.600 0.600 64.400 60.210 ;
        RECT  0.600 0.600 1.210 135.520 ;
        RECT  0.600 91.020 64.400 135.520 ;
        RECT  4.080 91.020 60.940 135.690 ;
        LAYER M3 ;
        RECT  0.600 247.660 14.720 249.400 ;
        RECT  50.220 247.660 64.400 249.400 ;
        RECT  0.600 0.600 64.400 60.480 ;
        RECT  2.000 0.000 63.000 88.700 ;
        RECT  0.600 0.600 1.480 91.220 ;
        RECT  0.600 90.750 64.400 91.220 ;
        RECT  0.600 124.090 64.550 128.560 ;
        RECT  0.600 124.090 64.400 129.850 ;
        RECT  1.400 124.090 63.600 135.790 ;
        RECT  62.370 124.090 63.600 154.120 ;
        RECT  1.400 124.090 2.470 154.470 ;
        RECT  1.640 155.040 63.360 171.560 ;
        RECT  3.070 124.090 58.100 185.950 ;
        RECT  1.640 183.580 63.360 185.950 ;
        RECT  3.070 124.090 5.960 195.660 ;
        RECT  10.490 144.980 61.290 200.820 ;
        RECT  1.640 196.170 63.360 200.820 ;
        RECT  58.010 144.980 59.020 201.060 ;
        RECT  60.060 144.980 61.290 201.060 ;
        LAYER TOP_M ;
        RECT  2.970 247.550 14.690 249.400 ;
        RECT  0.600 247.690 14.690 249.400 ;
        RECT  2.970 222.720 62.030 246.820 ;
        RECT  2.970 201.660 62.030 221.520 ;
        RECT  2.970 123.850 62.030 200.930 ;
        RECT  2.970 92.060 62.030 123.250 ;
        RECT  50.250 247.550 62.030 249.400 ;
        RECT  50.250 247.690 64.400 249.400 ;
        RECT  2.000 0.000 63.000 91.190 ;
        RECT  0.600 0.600 64.400 91.190 ;
        RECT  2.970 0.000 62.030 91.330 ;
    END
END pvdc

MACRO pvda
    CLASS PAD ;
    FOREIGN pvda 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 65.000 BY 250.000 ;
    SYMMETRY X Y R90 ;
    SITE IOSite_c ;
    PIN VDDO
        DIRECTION OUTPUT ;
        USE power ;
        PORT
        LAYER M3 ;
        RECT  64.200 192.330 65.000 200.640 ;
        RECT  0.000 201.660 65.000 221.520 ;
        RECT  0.000 222.720 65.000 246.820 ;
        RECT  0.000 192.330 0.800 200.640 ;
        LAYER M2 ;
        RECT  0.000 186.470 65.000 195.650 ;
        RECT  2.000 61.000 63.000 90.230 ;
        LAYER TOP_M ;
        RECT  0.000 195.170 65.000 200.640 ;
        RECT  0.000 201.660 65.000 221.520 ;
        RECT  0.000 222.720 65.000 246.820 ;
        END
    END VDDO
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        PORT
        LAYER M3 ;
        RECT  64.200 163.510 65.000 190.890 ;
        RECT  0.000 163.510 0.800 190.890 ;
        LAYER M2 ;
        RECT  0.000 172.080 65.000 183.060 ;
        LAYER TOP_M ;
        RECT  0.000 163.500 65.000 194.560 ;
        END
    END VDD
    PIN VSSO
        DIRECTION INOUT ;
        USE ground ;
        PORT
        LAYER M3 ;
        RECT  64.200 92.060 65.000 123.250 ;
        RECT  0.000 92.060 65.000 122.850 ;
        RECT  0.000 92.060 2.470 123.250 ;
        RECT  64.200 149.940 65.000 162.610 ;
        RECT  0.000 149.940 0.800 162.610 ;
        LAYER M2 ;
        RECT  0.000 147.040 65.000 154.520 ;
        LAYER TOP_M ;
        RECT  0.000 92.060 65.000 123.250 ;
        RECT  0.000 155.410 65.000 162.610 ;
        END
    END VSSO
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        PORT
        LAYER M3 ;
        RECT  64.200 130.690 65.000 148.880 ;
        RECT  0.000 130.690 0.800 148.880 ;
        LAYER M2 ;
        RECT  0.000 136.310 65.000 146.340 ;
        LAYER TOP_M ;
        RECT  0.000 123.850 65.000 154.560 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  2.000 0.000 63.000 250.000 ;
        RECT  0.000 88.990 65.000 130.360 ;
        RECT  0.000 136.510 65.000 157.550 ;
        RECT  0.500 136.510 64.500 163.550 ;
        RECT  0.600 0.600 64.400 250.000 ;
        RECT  0.000 198.470 65.000 250.000 ;
        LAYER M2 ;
        RECT  7.270 196.250 9.370 249.400 ;
        RECT  55.630 196.250 57.730 249.400 ;
        RECT  0.600 196.440 64.400 249.400 ;
        RECT  0.600 183.850 64.400 185.680 ;
        RECT  0.600 155.310 64.400 171.290 ;
        RECT  2.000 0.000 63.000 60.210 ;
        RECT  0.600 0.600 64.400 60.210 ;
        RECT  0.600 0.600 1.210 135.520 ;
        RECT  0.600 91.020 64.400 135.520 ;
        RECT  4.080 91.020 60.940 135.690 ;
        LAYER M3 ;
        RECT  0.600 247.660 64.400 249.400 ;
        RECT  0.600 124.090 64.400 129.850 ;
        RECT  3.310 123.690 63.360 135.790 ;
        RECT  1.400 124.090 63.360 135.790 ;
        RECT  1.400 124.090 2.470 154.470 ;
        RECT  1.640 155.040 63.360 171.560 ;
        RECT  1.640 183.580 63.360 185.950 ;
        RECT  3.110 124.090 63.160 200.820 ;
        RECT  1.640 196.170 63.360 200.820 ;
        RECT  55.630 123.690 57.530 201.060 ;
        RECT  58.010 123.690 59.020 201.060 ;
        RECT  60.060 123.690 61.290 201.060 ;
        RECT  0.600 0.600 64.400 60.480 ;
        RECT  2.000 0.000 63.000 88.700 ;
        RECT  0.600 0.600 1.480 91.220 ;
        RECT  0.600 90.750 64.400 91.220 ;
        LAYER TOP_M ;
        RECT  0.600 247.690 64.400 249.400 ;
        RECT  2.000 0.000 63.000 91.190 ;
        RECT  0.600 0.600 64.400 91.190 ;
    END
END pvda

MACRO pvcf
    CLASS PAD ;
    FOREIGN pvcf 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.060 BY 250.000 ;
    SYMMETRY X Y R90 ;
    SITE IOSite_c ;
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        PORT
        LAYER M2 ;
        RECT  0.000 136.310 5.060 146.340 ;
        LAYER M3 ;
        RECT  0.000 130.690 5.060 148.880 ;
        LAYER TOP_M ;
        RECT  0.000 123.850 5.060 154.560 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  -0.470 88.990 5.530 130.360 ;
        RECT  0.600 0.600 4.460 250.000 ;
        RECT  -0.470 198.470 5.530 250.000 ;
        LAYER M2 ;
        RECT  0.600 147.130 4.460 249.400 ;
        RECT  0.600 0.600 4.460 135.520 ;
        LAYER M3 ;
        RECT  0.600 149.720 4.460 249.400 ;
        RECT  0.600 0.600 4.460 129.850 ;
        LAYER TOP_M ;
        RECT  0.600 155.430 4.460 249.400 ;
        RECT  0.600 0.600 4.460 122.980 ;
    END
END pvcf

MACRO pvce
    CLASS PAD ;
    FOREIGN pvce 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.060 BY 250.000 ;
    SYMMETRY X Y R90 ;
    SITE IOSite_c ;
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        PORT
        LAYER M2 ;
        RECT  0.000 136.310 5.060 146.340 ;
        LAYER M3 ;
        RECT  0.000 130.690 5.060 148.880 ;
        LAYER TOP_M ;
        RECT  0.000 123.850 5.060 154.560 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        PORT
        LAYER M2 ;
        RECT  0.000 172.080 5.060 183.060 ;
        LAYER M3 ;
        RECT  0.000 163.510 5.060 190.890 ;
        LAYER TOP_M ;
        RECT  0.000 163.500 5.060 194.560 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  -0.470 88.990 5.530 130.360 ;
        RECT  0.600 0.600 4.460 250.000 ;
        RECT  -0.470 198.470 5.530 250.000 ;
        LAYER M2 ;
        RECT  0.600 183.850 4.460 249.400 ;
        RECT  0.600 147.130 4.460 171.290 ;
        RECT  0.600 0.600 4.460 135.520 ;
        LAYER M3 ;
        RECT  0.600 191.730 4.460 249.400 ;
        RECT  0.600 149.720 4.460 162.670 ;
        RECT  0.600 0.600 4.460 129.850 ;
        LAYER TOP_M ;
        RECT  0.600 195.430 4.460 249.400 ;
        RECT  0.600 155.430 4.460 162.630 ;
        RECT  0.600 0.600 4.460 122.980 ;
    END
END pvce

MACRO pv0i
    CLASS PAD ;
    FOREIGN pv0i 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 65.000 BY 250.000 ;
    SYMMETRY X Y R90 ;
    SITE IOSite_c ;
    PIN VDDO
        DIRECTION INOUT ;
        USE power ;
        PORT
        LAYER M3 ;
        RECT  64.200 192.330 65.000 200.640 ;
        RECT  0.000 201.660 65.000 221.520 ;
        RECT  0.000 222.720 65.000 246.820 ;
        RECT  0.000 192.330 0.800 200.640 ;
        LAYER M2 ;
        RECT  0.000 186.470 65.000 195.650 ;
        LAYER TOP_M ;
        RECT  0.000 195.170 65.000 200.640 ;
        RECT  0.000 201.660 65.000 221.520 ;
        RECT  0.000 222.720 65.000 246.820 ;
        END
    END VDDO
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        PORT
        LAYER M3 ;
        RECT  64.200 163.510 65.000 190.890 ;
        RECT  0.000 163.510 3.220 190.890 ;
        LAYER M2 ;
        RECT  0.000 172.080 65.000 183.060 ;
        LAYER TOP_M ;
        RECT  0.000 163.500 65.000 194.560 ;
        END
    END VDD
    PIN VSSO
        DIRECTION INOUT ;
        USE ground ;
        PORT
        LAYER M3 ;
        RECT  64.200 92.060 65.000 123.250 ;
        RECT  0.000 92.060 65.000 117.850 ;
        RECT  0.000 92.060 2.470 123.250 ;
        RECT  64.200 149.940 65.000 162.610 ;
        RECT  0.000 149.940 0.800 162.610 ;
        LAYER M2 ;
        RECT  0.000 147.040 65.000 154.520 ;
        LAYER TOP_M ;
        RECT  0.000 92.060 65.000 123.250 ;
        RECT  0.000 155.410 65.000 162.610 ;
        END
    END VSSO
    PIN VSS
        DIRECTION OUTPUT ;
        USE ground ;
        PORT
	CLASS CORE ;
        LAYER M3 ;
        RECT  64.200 130.690 65.000 148.880 ;
        RECT  15.560 247.420 49.380 250.000 ;
        RECT  0.000 130.690 0.800 148.880 ;
        LAYER M2 ;
        RECT  0.000 136.310 65.000 146.340 ;
        RECT  2.000 61.000 63.000 90.230 ;
        RECT  15.560 246.630 49.380 250.000 ;
        LAYER TOP_M ;
        RECT  0.000 123.850 65.000 154.560 ;
        RECT  15.560 247.420 49.380 250.000 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  2.000 0.000 63.000 250.000 ;
        RECT  0.000 88.990 65.000 130.360 ;
        RECT  0.000 136.510 65.000 157.550 ;
        RECT  0.500 136.510 64.500 163.550 ;
        RECT  0.600 0.600 64.400 250.000 ;
        RECT  0.000 198.470 65.000 250.000 ;
        LAYER M2 ;
        RECT  5.280 196.250 9.830 249.400 ;
        RECT  0.600 196.440 64.400 245.840 ;
        RECT  0.600 196.440 14.950 246.720 ;
        RECT  50.060 196.440 64.400 246.720 ;
        RECT  0.600 196.440 14.770 249.400 ;
        RECT  50.170 196.440 64.400 249.400 ;
        RECT  0.600 183.850 64.400 185.680 ;
        RECT  0.600 155.310 64.400 171.290 ;
        RECT  2.000 0.000 63.000 60.210 ;
        RECT  0.600 0.600 64.400 60.210 ;
        RECT  0.600 0.600 1.210 135.520 ;
        RECT  0.600 91.020 64.400 135.520 ;
        RECT  1.540 91.020 63.110 135.690 ;
        LAYER M3 ;
        RECT  0.600 247.660 14.720 249.400 ;
        RECT  50.220 247.660 64.400 249.400 ;
        RECT  0.600 124.090 64.400 129.850 ;
        RECT  3.070 118.690 63.360 135.790 ;
        RECT  1.400 124.090 63.360 135.790 ;
        RECT  1.400 124.090 2.470 154.470 ;
        RECT  3.070 118.510 62.880 162.670 ;
        RECT  1.640 155.040 63.360 162.670 ;
        RECT  4.060 155.040 63.360 182.880 ;
        RECT  4.060 118.510 56.875 200.820 ;
        RECT  4.060 183.580 63.360 185.950 ;
        RECT  4.060 183.580 60.010 200.820 ;
        RECT  3.070 191.730 60.010 200.820 ;
        RECT  1.640 196.170 63.360 200.820 ;
        RECT  58.930 183.580 60.010 201.060 ;
        RECT  0.600 0.600 64.400 60.480 ;
        RECT  2.000 0.000 63.000 88.700 ;
        RECT  0.600 0.600 1.480 91.220 ;
        RECT  0.600 90.750 64.400 91.220 ;
        LAYER TOP_M ;
        RECT  0.600 247.690 14.690 249.400 ;
        RECT  50.250 247.690 64.400 249.400 ;
        RECT  2.000 0.000 63.000 91.190 ;
        RECT  0.600 0.600 64.400 91.190 ;
    END
END pv0i

MACRO pv0f
    CLASS PAD ;
    FOREIGN pv0f 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 65.000 BY 250.000 ;
    SYMMETRY X Y R90 ;
    SITE IOSite_c ;
    PIN VDDO
        DIRECTION INOUT ;
        USE power ;
        PORT
        LAYER M3 ;
        RECT  64.200 192.330 65.000 200.640 ;
        RECT  0.000 201.660 65.000 221.520 ;
        RECT  0.000 222.720 65.000 246.820 ;
        RECT  0.000 192.330 0.800 200.640 ;
        LAYER M2 ;
        RECT  0.000 186.470 65.000 195.650 ;
        LAYER TOP_M ;
        RECT  0.000 195.170 65.000 200.640 ;
        RECT  0.000 201.660 65.000 221.520 ;
        RECT  0.000 222.720 65.000 246.820 ;
        END
    END VDDO
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        PORT
        LAYER M3 ;
        RECT  64.200 163.510 65.000 190.890 ;
        RECT  0.000 163.510 0.800 190.890 ;
        LAYER M2 ;
        RECT  0.000 172.080 65.000 183.060 ;
        LAYER TOP_M ;
        RECT  0.000 163.500 65.000 194.560 ;
        END
    END VDD
    PIN VSS
        DIRECTION OUTPUT ;
        USE ground ;
        PORT
        LAYER M3 ;
        RECT  64.200 92.060 65.000 123.250 ;
        RECT  0.000 92.060 65.000 117.850 ;
        RECT  0.000 92.060 2.470 123.250 ;
        RECT  64.200 130.690 65.000 148.880 ;
        RECT  64.200 149.940 65.000 162.610 ;
        RECT  0.000 130.690 0.800 148.880 ;
        RECT  0.000 149.940 0.800 162.610 ;
        LAYER M2 ;
        RECT  0.000 136.310 65.000 146.340 ;
        RECT  0.000 147.040 65.000 154.520 ;
        RECT  2.000 61.000 63.000 90.230 ;
        LAYER TOP_M ;
        RECT  0.000 92.060 65.000 123.250 ;
        RECT  0.000 123.850 65.000 154.560 ;
        RECT  0.000 155.410 65.000 162.610 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  2.000 0.000 63.000 250.000 ;
        RECT  0.000 88.990 65.000 130.360 ;
        RECT  0.000 136.510 65.000 157.550 ;
        RECT  0.500 136.510 64.500 163.550 ;
        RECT  0.600 0.600 64.400 250.000 ;
        RECT  0.000 198.470 65.000 250.000 ;
        LAYER M2 ;
        RECT  0.600 196.440 64.400 249.400 ;
        RECT  0.600 183.850 64.400 185.680 ;
        RECT  0.600 155.310 64.400 171.290 ;
        RECT  2.000 0.000 63.000 60.210 ;
        RECT  0.600 0.600 64.400 60.210 ;
        RECT  0.600 0.600 1.210 135.520 ;
        RECT  0.600 91.020 64.400 135.520 ;
        LAYER M3 ;
        RECT  0.600 247.660 64.400 249.400 ;
        RECT  0.600 124.090 64.400 129.850 ;
        RECT  1.400 124.090 63.520 135.790 ;
        RECT  1.400 124.090 2.470 154.470 ;
        RECT  1.640 155.040 63.520 171.560 ;
        RECT  1.640 183.580 63.520 185.950 ;
        RECT  3.300 124.090 63.520 200.820 ;
        RECT  3.310 118.640 63.520 200.820 ;
        RECT  1.640 196.170 63.520 200.820 ;
        RECT  55.270 118.640 56.355 201.060 ;
        RECT  0.600 0.600 64.400 60.480 ;
        RECT  2.000 0.000 63.000 88.700 ;
        RECT  0.600 0.600 1.480 91.220 ;
        RECT  0.600 90.750 64.400 91.220 ;
        LAYER TOP_M ;
        RECT  0.600 247.690 64.400 249.400 ;
        RECT  2.000 0.000 63.000 91.190 ;
        RECT  0.600 0.600 64.400 91.190 ;
    END
END pv0f

MACRO pv0c
    CLASS PAD ;
    FOREIGN pv0c 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 65.000 BY 250.000 ;
    SYMMETRY X Y R90 ;
    SITE IOSite_c ;
    PIN VDDO
        DIRECTION INOUT ;
        USE power ;
        PORT
        LAYER M3 ;
        RECT  64.200 192.330 65.000 200.640 ;
        RECT  0.000 201.660 65.000 221.520 ;
        RECT  0.000 222.720 65.000 246.820 ;
        RECT  0.000 192.330 0.800 200.640 ;
        LAYER M2 ;
        RECT  0.000 186.470 65.000 195.650 ;
        LAYER TOP_M ;
        RECT  0.000 195.170 65.000 200.640 ;
        RECT  0.000 201.660 65.000 221.520 ;
        RECT  0.000 222.720 65.000 246.820 ;
        END
    END VDDO
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        PORT
        LAYER M3 ;
        RECT  64.200 163.510 65.000 190.890 ;
        RECT  0.000 163.510 3.110 190.890 ;
        LAYER M2 ;
        RECT  0.000 172.080 65.000 183.060 ;
        LAYER TOP_M ;
        RECT  0.000 163.500 65.000 194.560 ;
        END
    END VDD
    PIN VSSO
        DIRECTION INOUT ;
        USE ground ;
        PORT
        LAYER M3 ;
        RECT  64.200 92.060 65.000 123.250 ;
        RECT  0.000 92.060 65.000 117.850 ;
        RECT  0.000 92.060 2.470 123.250 ;
        RECT  64.200 149.940 65.000 162.610 ;
        RECT  0.000 149.940 0.800 162.610 ;
        LAYER M2 ;
        RECT  57.230 147.040 65.000 154.520 ;
        RECT  0.000 147.040 65.000 149.960 ;
        RECT  0.000 147.040 7.630 154.520 ;
        LAYER TOP_M ;
        RECT  0.000 92.060 65.000 123.250 ;
        RECT  0.000 155.410 65.000 162.610 ;
        END
    END VSSO
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        PORT
        LAYER M3 ;
        RECT  64.200 130.690 65.000 148.880 ;
        RECT  0.000 130.690 0.800 148.880 ;
        LAYER M2 ;
        RECT  0.000 136.310 65.000 146.340 ;
        LAYER TOP_M ;
        RECT  0.000 123.850 65.000 154.560 ;
        END
    END VSS
    PIN VSSC
        DIRECTION OUTPUT ;
        USE ground ;
        PORT
	CLASS CORE ;
        LAYER M3 ;
        RECT  15.560 247.420 49.380 250.000 ;
        LAYER M2 ;
        RECT  2.000 61.000 63.000 90.230 ;
        RECT  15.560 246.630 49.380 250.000 ;
        LAYER TOP_M ;
        RECT  15.560 247.420 49.380 250.000 ;
        END
    END VSSC
    OBS
        LAYER M1 ;
        RECT  2.000 0.000 63.000 250.000 ;
        RECT  0.000 88.990 65.000 130.360 ;
        RECT  0.000 136.510 65.000 157.550 ;
        RECT  0.500 136.510 64.500 163.550 ;
        RECT  0.600 0.600 64.400 250.000 ;
        RECT  0.000 198.470 65.000 250.000 ;
        LAYER M2 ;
        RECT  5.280 196.250 9.830 249.400 ;
        RECT  55.030 196.250 56.930 249.400 ;
        RECT  0.600 196.440 64.400 245.840 ;
        RECT  0.600 196.440 14.950 246.720 ;
        RECT  50.060 196.440 64.400 246.720 ;
        RECT  0.600 196.440 14.770 249.400 ;
        RECT  50.170 196.440 64.400 249.400 ;
        RECT  0.600 183.850 64.400 185.680 ;
        RECT  8.230 150.560 56.630 154.520 ;
        RECT  8.420 150.560 56.440 171.290 ;
        RECT  0.600 155.310 64.400 171.290 ;
        RECT  2.000 0.000 63.000 60.210 ;
        RECT  0.600 0.600 64.400 60.210 ;
        RECT  0.600 0.600 1.210 135.520 ;
        RECT  0.600 91.020 64.400 135.520 ;
        RECT  1.540 91.020 63.110 135.690 ;
        LAYER M3 ;
        RECT  0.600 247.660 14.720 249.400 ;
        RECT  50.220 247.660 64.400 249.400 ;
        RECT  0.600 124.090 64.400 129.850 ;
        RECT  3.070 118.690 63.360 135.790 ;
        RECT  1.400 124.090 63.360 135.790 ;
        RECT  1.400 124.090 2.470 154.470 ;
        RECT  3.070 118.510 62.880 162.670 ;
        RECT  1.640 155.040 63.360 162.670 ;
        RECT  3.950 155.040 63.360 182.880 ;
        RECT  3.950 118.510 56.880 200.820 ;
        RECT  3.950 183.580 63.360 185.950 ;
        RECT  3.950 183.580 60.010 200.820 ;
        RECT  3.070 191.730 60.010 200.820 ;
        RECT  1.640 196.170 63.360 200.820 ;
        RECT  58.930 183.580 60.010 201.060 ;
        RECT  0.600 0.600 64.400 60.480 ;
        RECT  2.000 0.000 63.000 88.700 ;
        RECT  0.600 0.600 1.480 91.220 ;
        RECT  0.600 90.750 64.400 91.220 ;
        LAYER TOP_M ;
        RECT  0.600 247.690 14.690 249.400 ;
        RECT  50.250 247.690 64.400 249.400 ;
        RECT  2.000 0.000 63.000 91.190 ;
        RECT  0.600 0.600 64.400 91.190 ;
    END
END pv0c

MACRO pv0a
    CLASS PAD ;
    FOREIGN pv0a 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 65.000 BY 250.000 ;
    SYMMETRY X Y R90 ;
    SITE IOSite_c ;
    PIN VDDO
        DIRECTION INOUT ;
        USE power ;
        PORT
        LAYER M3 ;
        RECT  64.200 192.330 65.000 200.640 ;
        RECT  0.000 201.660 65.000 221.520 ;
        RECT  0.000 222.720 65.000 246.820 ;
        RECT  0.000 192.330 0.800 200.640 ;
        LAYER M2 ;
        RECT  0.000 186.470 65.000 195.650 ;
        LAYER TOP_M ;
        RECT  0.000 195.170 65.000 200.640 ;
        RECT  0.000 201.660 65.000 221.520 ;
        RECT  0.000 222.720 65.000 246.820 ;
        END
    END VDDO
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        PORT
        LAYER M3 ;
        RECT  64.200 163.510 65.000 190.890 ;
        RECT  0.000 163.510 0.800 190.890 ;
        LAYER M2 ;
        RECT  0.000 172.080 65.000 183.060 ;
        LAYER TOP_M ;
        RECT  0.000 163.500 65.000 194.560 ;
        END
    END VDD
    PIN VSSO
        DIRECTION OUTPUT ;
        USE ground ;
        PORT
        LAYER M3 ;
        RECT  64.200 92.060 65.000 123.250 ;
        RECT  0.000 92.060 65.000 117.850 ;
        RECT  0.000 92.060 2.470 123.250 ;
        RECT  64.200 149.940 65.000 162.610 ;
        RECT  0.000 149.940 0.800 162.610 ;
        LAYER M2 ;
        RECT  0.000 147.040 65.000 154.520 ;
        RECT  2.000 61.000 63.000 90.230 ;
        LAYER TOP_M ;
        RECT  0.000 92.060 65.000 123.250 ;
        RECT  0.000 155.410 65.000 162.610 ;
        END
    END VSSO
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        PORT
        LAYER M3 ;
        RECT  64.200 130.690 65.000 148.880 ;
        RECT  0.000 130.690 0.800 148.880 ;
        LAYER M2 ;
        RECT  0.000 136.310 65.000 146.340 ;
        LAYER TOP_M ;
        RECT  0.000 123.850 65.000 154.560 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  2.000 0.000 63.000 250.000 ;
        RECT  0.000 88.990 65.000 130.360 ;
        RECT  0.000 136.510 65.000 157.550 ;
        RECT  0.500 136.510 64.500 163.550 ;
        RECT  0.600 0.600 64.400 250.000 ;
        RECT  0.000 198.470 65.000 250.000 ;
        LAYER M2 ;
        RECT  0.600 196.440 64.400 249.400 ;
        RECT  0.600 183.850 64.400 185.680 ;
        RECT  0.600 155.310 64.400 171.290 ;
        RECT  2.000 0.000 63.000 60.210 ;
        RECT  0.600 0.600 64.400 60.210 ;
        RECT  0.600 0.600 1.210 135.520 ;
        RECT  0.600 91.020 64.400 135.520 ;
        RECT  2.560 91.020 62.460 135.690 ;
        LAYER M3 ;
        RECT  0.600 247.660 64.400 249.400 ;
        RECT  0.600 124.090 64.400 129.850 ;
        RECT  1.400 124.090 63.455 135.790 ;
        RECT  1.400 124.090 2.470 154.470 ;
        RECT  1.640 155.040 63.455 171.560 ;
        RECT  1.640 183.580 63.455 185.950 ;
        RECT  3.300 124.090 63.455 200.820 ;
        RECT  3.310 118.450 63.455 200.820 ;
        RECT  1.640 196.170 63.455 200.820 ;
        RECT  55.270 118.450 56.355 201.060 ;
        RECT  0.600 0.600 64.400 60.480 ;
        RECT  2.000 0.000 63.000 88.700 ;
        RECT  0.600 0.600 1.480 91.220 ;
        RECT  0.600 90.750 64.400 91.220 ;
        LAYER TOP_M ;
        RECT  0.600 247.690 64.400 249.400 ;
        RECT  2.000 0.000 63.000 91.190 ;
        RECT  0.600 0.600 64.400 91.190 ;
    END
END pv0a

MACRO pt3t03u
    CLASS PAD ;
    FOREIGN pt3t03u 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 65.000 BY 250.000 ;
    SYMMETRY X Y R90 ;
    SITE IOSite_c ;
    PIN PAD
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 55.440  LAYER TOP_M  ;
        ANTENNAPARTIALMETALSIDEAREA 287.938  LAYER M3  ;
        ANTENNAPARTIALMETALSIDEAREA 480.740  LAYER M2  ;
        ANTENNADIFFAREA 2657.280  LAYER TOP_M  ;
        ANTENNADIFFAREA 2657.280  LAYER M3  ;
        ANTENNADIFFAREA 1209.600  LAYER M2  ;
        ANTENNAPARTIALCUTAREA 632.318  LAYER TOP_V  ;
        ANTENNAPARTIALCUTAREA 349.898  LAYER V3  ;
        ANTENNAPARTIALCUTAREA 255.798  LAYER V2  ;
        PORT
        LAYER M3 ;
        RECT  23.740 249.580 25.740 250.000 ;
        LAYER M2 ;
        RECT  2.000 61.000 63.000 90.230 ;
        RECT  23.740 246.275 25.740 250.000 ;
        END
    END PAD
    PIN OEN
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 81.726  LAYER M2  ;
        ANTENNAPARTIALMETALSIDEAREA 67.374  LAYER M1  ;
        ANTENNAPARTIALMETALSIDEAREA 41.679  LAYER M3  ;
        ANTENNADIFFAREA 0.250  LAYER M3  ;
        ANTENNAPARTIALCUTAREA 0.135  LAYER V3  ;
        ANTENNAPARTIALCUTAREA 0.203  LAYER V2  ;
        ANTENNAGATEAREA 8.100  LAYER M2  ;
        ANTENNAGATEAREA 9.900  LAYER M3  ;
        PORT
        LAYER M3 ;
        RECT  28.870 249.580 29.600 250.000 ;
        LAYER M2 ;
        RECT  28.870 249.580 29.600 250.000 ;
        END
    END OEN
    PIN I
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 67.374  LAYER M1  ;
        ANTENNAPARTIALMETALSIDEAREA 80.804  LAYER M2  ;
        ANTENNAPARTIALMETALSIDEAREA 41.096  LAYER M3  ;
        ANTENNADIFFAREA 0.250  LAYER M3  ;
        ANTENNAPARTIALCUTAREA 0.270  LAYER V2  ;
        ANTENNAPARTIALCUTAREA 0.135  LAYER V3  ;
        ANTENNAGATEAREA 18.900  LAYER M2  ;
        ANTENNAGATEAREA 20.700  LAYER M3  ;
        PORT
        LAYER M3 ;
        RECT  27.840 249.580 28.570 250.000 ;
        LAYER M2 ;
        RECT  27.840 249.580 28.570 250.000 ;
        END
    END I
    PIN VDDO
        DIRECTION INOUT ;
        USE power ;
        PORT
        LAYER M3 ;
        RECT  64.200 192.330 65.000 200.640 ;
        RECT  0.000 201.660 65.000 221.520 ;
        RECT  0.000 222.720 65.000 246.820 ;
        RECT  0.000 192.330 0.800 200.640 ;
        LAYER M2 ;
        RECT  0.000 186.470 65.000 195.650 ;
        LAYER TOP_M ;
        RECT  0.000 195.170 65.000 200.640 ;
        RECT  0.000 201.660 65.000 221.520 ;
        RECT  0.000 222.720 65.000 246.820 ;
        END
    END VDDO
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        PORT
        LAYER M3 ;
        RECT  64.200 163.510 65.000 190.890 ;
        RECT  0.000 163.510 0.800 190.890 ;
        LAYER M2 ;
        RECT  0.000 172.080 65.000 183.060 ;
        LAYER TOP_M ;
        RECT  0.000 163.500 65.000 194.560 ;
        END
    END VDD
    PIN VSSO
        DIRECTION INOUT ;
        USE ground ;
        PORT
        LAYER M3 ;
        RECT  0.000 92.060 65.000 123.250 ;
        RECT  64.200 149.940 65.000 162.610 ;
        RECT  0.000 149.940 0.800 162.610 ;
        LAYER M2 ;
        RECT  0.000 147.040 65.000 154.520 ;
        LAYER TOP_M ;
        RECT  0.000 92.060 65.000 123.250 ;
        RECT  0.000 155.410 65.000 162.610 ;
        END
    END VSSO
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        PORT
        LAYER M3 ;
        RECT  64.200 130.690 65.000 148.880 ;
        RECT  0.000 130.690 0.800 148.880 ;
        LAYER M2 ;
        RECT  0.000 136.310 65.000 146.340 ;
        LAYER TOP_M ;
        RECT  0.000 123.850 65.000 154.560 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  2.000 0.000 63.000 250.000 ;
        RECT  0.000 88.990 65.000 130.360 ;
        RECT  0.000 136.510 65.000 157.550 ;
        RECT  0.315 158.150 64.700 158.460 ;
        RECT  0.300 158.930 64.700 159.230 ;
        RECT  0.300 159.530 64.700 159.830 ;
        RECT  0.300 160.130 64.700 160.430 ;
        RECT  0.300 160.730 64.700 161.030 ;
        RECT  0.300 161.330 64.700 161.630 ;
        RECT  0.300 161.910 64.700 162.190 ;
        RECT  0.300 162.490 64.700 162.770 ;
        RECT  0.300 163.070 64.700 163.350 ;
        RECT  0.300 163.650 64.700 163.950 ;
        RECT  0.300 164.250 64.700 164.550 ;
        RECT  0.300 164.850 64.700 165.150 ;
        RECT  0.300 165.450 64.700 165.750 ;
        RECT  0.300 166.050 64.700 166.350 ;
        RECT  0.300 166.650 64.700 166.960 ;
        RECT  0.300 167.260 64.700 167.560 ;
        RECT  0.300 167.860 64.700 168.160 ;
        RECT  0.000 169.150 65.000 197.240 ;
        RECT  0.600 0.600 64.400 250.000 ;
        RECT  0.000 198.470 65.000 250.000 ;
        LAYER M2 ;
        RECT  63.180 196.430 63.670 249.400 ;
        RECT  0.600 196.440 64.400 245.485 ;
        RECT  26.530 196.440 64.400 248.790 ;
        RECT  0.600 196.440 22.950 249.400 ;
        RECT  26.530 196.440 27.050 249.400 ;
        RECT  30.390 196.440 64.400 249.400 ;
        RECT  0.600 183.850 64.400 185.680 ;
        RECT  46.230 183.850 51.730 185.870 ;
        RECT  4.480 154.920 7.530 171.290 ;
        RECT  8.170 155.125 8.490 171.290 ;
        RECT  21.210 155.160 21.560 171.290 ;
        RECT  21.860 155.140 22.180 171.290 ;
        RECT  31.895 155.120 35.765 171.290 ;
        RECT  53.655 155.035 53.935 171.290 ;
        RECT  56.365 155.280 56.645 171.290 ;
        RECT  57.120 155.300 57.400 171.290 ;
        RECT  57.835 155.130 58.115 171.290 ;
        RECT  0.600 155.310 64.400 171.290 ;
        RECT  53.895 155.310 55.870 171.370 ;
        RECT  3.170 155.310 3.450 171.380 ;
        RECT  34.655 155.310 38.715 171.480 ;
        RECT  39.605 155.310 42.020 171.480 ;
        RECT  2.000 0.000 63.000 60.210 ;
        RECT  0.600 0.600 64.400 60.210 ;
        RECT  0.600 0.600 1.210 135.520 ;
        RECT  0.600 91.020 64.400 135.520 ;
        RECT  4.080 91.020 60.940 135.690 ;
        RECT  62.580 91.020 62.995 135.710 ;
        LAYER M3 ;
        RECT  0.600 247.660 23.220 248.740 ;
        RECT  0.600 247.660 22.900 249.400 ;
        RECT  26.260 247.660 64.400 248.740 ;
        RECT  26.580 247.660 27.000 249.400 ;
        RECT  30.440 247.660 64.400 249.400 ;
        RECT  0.600 124.090 64.400 129.850 ;
        RECT  1.640 124.090 63.600 135.790 ;
        RECT  1.810 124.090 2.830 154.520 ;
        RECT  3.510 124.090 63.600 171.560 ;
        RECT  4.040 123.970 60.900 171.560 ;
        RECT  1.640 155.040 63.600 171.560 ;
        RECT  1.640 183.580 63.600 185.950 ;
        RECT  5.515 124.090 63.600 200.820 ;
        RECT  1.640 196.170 63.600 200.820 ;
        RECT  0.600 0.600 64.400 60.480 ;
        RECT  2.000 0.000 63.000 88.700 ;
        RECT  0.600 0.600 1.480 91.220 ;
        RECT  0.600 90.750 64.400 91.220 ;
        LAYER TOP_M ;
        RECT  0.600 247.690 64.400 248.850 ;
        RECT  0.600 247.690 23.010 249.400 ;
        RECT  26.470 247.690 27.110 249.400 ;
        RECT  30.330 247.690 64.400 249.400 ;
        RECT  2.000 0.000 63.000 91.190 ;
        RECT  0.600 0.600 64.400 91.190 ;
    END
END pt3t03u

MACRO pt3t03d
    CLASS PAD ;
    FOREIGN pt3t03d 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 65.000 BY 250.000 ;
    SYMMETRY X Y R90 ;
    SITE IOSite_c ;
    PIN PAD
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 55.440  LAYER TOP_M  ;
        ANTENNAPARTIALMETALSIDEAREA 287.938  LAYER M3  ;
        ANTENNAPARTIALMETALSIDEAREA 480.740  LAYER M2  ;
        ANTENNADIFFAREA 2657.280  LAYER TOP_M  ;
        ANTENNADIFFAREA 2657.280  LAYER M3  ;
        ANTENNADIFFAREA 1209.600  LAYER M2  ;
        ANTENNAPARTIALCUTAREA 632.318  LAYER TOP_V  ;
        ANTENNAPARTIALCUTAREA 349.898  LAYER V3  ;
        ANTENNAPARTIALCUTAREA 255.798  LAYER V2  ;
        PORT
        LAYER M3 ;
        RECT  23.740 249.580 25.740 250.000 ;
        LAYER M2 ;
        RECT  2.000 61.000 63.000 90.230 ;
        RECT  23.740 246.275 25.740 250.000 ;
        END
    END PAD
    PIN OEN
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 81.726  LAYER M2  ;
        ANTENNAPARTIALMETALSIDEAREA 67.374  LAYER M1  ;
        ANTENNAPARTIALMETALSIDEAREA 41.679  LAYER M3  ;
        ANTENNADIFFAREA 0.250  LAYER M3  ;
        ANTENNAPARTIALCUTAREA 0.135  LAYER V3  ;
        ANTENNAPARTIALCUTAREA 0.203  LAYER V2  ;
        ANTENNAGATEAREA 8.100  LAYER M2  ;
        ANTENNAGATEAREA 9.900  LAYER M3  ;
        PORT
        LAYER M3 ;
        RECT  28.870 249.580 29.600 250.000 ;
        LAYER M2 ;
        RECT  28.870 249.580 29.600 250.000 ;
        END
    END OEN
    PIN I
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 67.374  LAYER M1  ;
        ANTENNAPARTIALMETALSIDEAREA 80.804  LAYER M2  ;
        ANTENNAPARTIALMETALSIDEAREA 41.096  LAYER M3  ;
        ANTENNADIFFAREA 0.250  LAYER M3  ;
        ANTENNAPARTIALCUTAREA 0.270  LAYER V2  ;
        ANTENNAPARTIALCUTAREA 0.135  LAYER V3  ;
        ANTENNAGATEAREA 18.900  LAYER M2  ;
        ANTENNAGATEAREA 20.700  LAYER M3  ;
        PORT
        LAYER M3 ;
        RECT  27.840 249.580 28.570 250.000 ;
        LAYER M2 ;
        RECT  27.840 249.580 28.570 250.000 ;
        END
    END I
    PIN VDDO
        DIRECTION INOUT ;
        USE power ;
        PORT
        LAYER M3 ;
        RECT  64.200 192.330 65.000 200.640 ;
        RECT  0.000 201.660 65.000 221.520 ;
        RECT  0.000 222.720 65.000 246.820 ;
        RECT  0.000 192.330 0.800 200.640 ;
        LAYER M2 ;
        RECT  0.000 186.470 65.000 195.650 ;
        LAYER TOP_M ;
        RECT  0.000 195.170 65.000 200.640 ;
        RECT  0.000 201.660 65.000 221.520 ;
        RECT  0.000 222.720 65.000 246.820 ;
        END
    END VDDO
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        PORT
        LAYER M3 ;
        RECT  64.200 163.510 65.000 190.890 ;
        RECT  0.000 163.510 0.800 190.890 ;
        LAYER M2 ;
        RECT  0.000 172.080 65.000 183.060 ;
        LAYER TOP_M ;
        RECT  0.000 163.500 65.000 194.560 ;
        END
    END VDD
    PIN VSSO
        DIRECTION INOUT ;
        USE ground ;
        PORT
        LAYER M3 ;
        RECT  0.000 92.060 65.000 123.250 ;
        RECT  64.200 149.940 65.000 162.610 ;
        RECT  0.000 149.940 0.800 162.610 ;
        LAYER M2 ;
        RECT  0.000 147.040 65.000 154.520 ;
        LAYER TOP_M ;
        RECT  0.000 92.060 65.000 123.250 ;
        RECT  0.000 155.410 65.000 162.610 ;
        END
    END VSSO
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        PORT
        LAYER M3 ;
        RECT  64.200 130.690 65.000 148.880 ;
        RECT  0.000 130.690 0.800 148.880 ;
        LAYER M2 ;
        RECT  0.000 136.310 65.000 146.340 ;
        LAYER TOP_M ;
        RECT  0.000 123.850 65.000 154.560 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  2.000 0.000 63.000 250.000 ;
        RECT  0.000 88.990 65.000 130.360 ;
        RECT  0.000 136.510 65.000 157.550 ;
        RECT  0.315 158.150 64.700 158.460 ;
        RECT  0.300 158.930 64.700 159.230 ;
        RECT  0.300 159.530 64.700 159.830 ;
        RECT  0.300 160.130 64.700 160.430 ;
        RECT  0.300 160.730 64.700 161.030 ;
        RECT  0.300 161.330 64.700 161.630 ;
        RECT  0.300 161.910 64.700 162.190 ;
        RECT  0.300 162.490 64.700 162.770 ;
        RECT  0.300 163.070 64.700 163.350 ;
        RECT  0.300 163.650 64.700 163.950 ;
        RECT  0.300 164.250 64.700 164.550 ;
        RECT  0.300 164.850 64.700 165.150 ;
        RECT  0.300 165.450 64.700 165.750 ;
        RECT  0.300 166.050 64.700 166.350 ;
        RECT  0.300 166.650 64.700 166.960 ;
        RECT  0.300 167.260 64.700 167.560 ;
        RECT  0.300 167.860 64.700 168.160 ;
        RECT  0.000 169.150 65.000 197.240 ;
        RECT  0.600 0.600 64.400 250.000 ;
        RECT  0.000 198.470 65.000 250.000 ;
        LAYER M2 ;
        RECT  63.180 196.430 63.670 249.400 ;
        RECT  0.600 196.440 64.400 245.485 ;
        RECT  26.530 196.440 64.400 248.790 ;
        RECT  0.600 196.440 22.950 249.400 ;
        RECT  26.530 196.440 27.050 249.400 ;
        RECT  30.390 196.440 64.400 249.400 ;
        RECT  0.600 183.850 64.400 185.680 ;
        RECT  46.230 183.850 51.730 185.870 ;
        RECT  4.480 154.920 7.530 171.290 ;
        RECT  8.170 155.125 8.490 171.290 ;
        RECT  21.210 155.160 21.560 171.290 ;
        RECT  21.860 155.140 22.180 171.290 ;
        RECT  31.895 155.120 35.765 171.290 ;
        RECT  49.255 155.125 51.495 171.290 ;
        RECT  52.435 155.295 52.745 171.290 ;
        RECT  53.655 155.035 53.935 171.290 ;
        RECT  56.365 155.280 56.645 171.290 ;
        RECT  57.120 155.300 57.400 171.290 ;
        RECT  57.835 155.130 58.115 171.290 ;
        RECT  0.600 155.310 64.400 171.290 ;
        RECT  53.895 155.310 55.870 171.370 ;
        RECT  3.170 155.310 3.450 171.380 ;
        RECT  34.655 155.310 38.715 171.480 ;
        RECT  39.605 155.310 42.020 171.480 ;
        RECT  2.000 0.000 63.000 60.210 ;
        RECT  0.600 0.600 64.400 60.210 ;
        RECT  0.600 0.600 1.210 135.520 ;
        RECT  0.600 91.020 64.400 135.520 ;
        RECT  4.080 91.020 60.940 135.690 ;
        RECT  62.580 91.020 62.995 135.710 ;
        LAYER M3 ;
        RECT  0.600 247.660 23.220 248.740 ;
        RECT  0.600 247.660 22.900 249.400 ;
        RECT  26.260 247.660 64.400 248.740 ;
        RECT  26.580 247.660 27.000 249.400 ;
        RECT  30.440 247.660 64.400 249.400 ;
        RECT  0.600 124.090 64.400 129.850 ;
        RECT  1.640 124.090 63.600 135.790 ;
        RECT  1.810 124.090 2.830 154.520 ;
        RECT  3.510 124.090 63.600 171.560 ;
        RECT  4.040 123.970 60.900 171.560 ;
        RECT  1.640 155.040 63.600 171.560 ;
        RECT  1.640 183.580 63.600 185.950 ;
        RECT  5.515 124.090 63.600 200.820 ;
        RECT  1.640 196.170 63.600 200.820 ;
        RECT  0.600 0.600 64.400 60.480 ;
        RECT  2.000 0.000 63.000 88.700 ;
        RECT  0.600 0.600 1.480 91.220 ;
        RECT  0.600 90.750 64.400 91.220 ;
        LAYER TOP_M ;
        RECT  0.600 247.690 64.400 248.850 ;
        RECT  0.600 247.690 23.010 249.400 ;
        RECT  26.470 247.690 27.110 249.400 ;
        RECT  30.330 247.690 64.400 249.400 ;
        RECT  2.000 0.000 63.000 91.190 ;
        RECT  0.600 0.600 64.400 91.190 ;
    END
END pt3t03d

MACRO pt3t03
    CLASS PAD ;
    FOREIGN pt3t03 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 65.000 BY 250.000 ;
    SYMMETRY X Y R90 ;
    SITE IOSite_c ;
    PIN PAD
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 55.440  LAYER TOP_M  ;
        ANTENNAPARTIALMETALSIDEAREA 287.938  LAYER M3  ;
        ANTENNAPARTIALMETALSIDEAREA 480.740  LAYER M2  ;
        ANTENNADIFFAREA 2657.280  LAYER TOP_M  ;
        ANTENNADIFFAREA 2657.280  LAYER M3  ;
        ANTENNADIFFAREA 1209.600  LAYER M2  ;
        ANTENNAPARTIALCUTAREA 632.318  LAYER TOP_V  ;
        ANTENNAPARTIALCUTAREA 349.898  LAYER V3  ;
        ANTENNAPARTIALCUTAREA 255.798  LAYER V2  ;
        PORT
        LAYER M3 ;
        RECT  23.740 249.580 25.740 250.000 ;
        LAYER M2 ;
        RECT  2.000 61.000 63.000 90.230 ;
        RECT  23.740 246.275 25.740 250.000 ;
        END
    END PAD
    PIN OEN
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 81.726  LAYER M2  ;
        ANTENNAPARTIALMETALSIDEAREA 67.374  LAYER M1  ;
        ANTENNAPARTIALMETALSIDEAREA 41.679  LAYER M3  ;
        ANTENNADIFFAREA 0.250  LAYER M3  ;
        ANTENNAPARTIALCUTAREA 0.135  LAYER V3  ;
        ANTENNAPARTIALCUTAREA 0.203  LAYER V2  ;
        ANTENNAGATEAREA 8.100  LAYER M2  ;
        ANTENNAGATEAREA 9.900  LAYER M3  ;
        PORT
        LAYER M3 ;
        RECT  28.870 249.580 29.600 250.000 ;
        LAYER M2 ;
        RECT  28.870 249.580 29.600 250.000 ;
        END
    END OEN
    PIN I
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 67.374  LAYER M1  ;
        ANTENNAPARTIALMETALSIDEAREA 80.804  LAYER M2  ;
        ANTENNAPARTIALMETALSIDEAREA 41.096  LAYER M3  ;
        ANTENNADIFFAREA 0.250  LAYER M3  ;
        ANTENNAPARTIALCUTAREA 0.270  LAYER V2  ;
        ANTENNAPARTIALCUTAREA 0.135  LAYER V3  ;
        ANTENNAGATEAREA 18.900  LAYER M2  ;
        ANTENNAGATEAREA 20.700  LAYER M3  ;
        PORT
        LAYER M3 ;
        RECT  27.840 249.580 28.570 250.000 ;
        LAYER M2 ;
        RECT  27.840 249.580 28.570 250.000 ;
        END
    END I
    PIN VDDO
        DIRECTION INOUT ;
        USE power ;
        PORT
        LAYER M3 ;
        RECT  64.200 192.330 65.000 200.640 ;
        RECT  0.000 201.660 65.000 221.520 ;
        RECT  0.000 222.720 65.000 246.820 ;
        RECT  0.000 192.330 0.800 200.640 ;
        LAYER M2 ;
        RECT  0.000 186.470 65.000 195.650 ;
        LAYER TOP_M ;
        RECT  0.000 195.170 65.000 200.640 ;
        RECT  0.000 201.660 65.000 221.520 ;
        RECT  0.000 222.720 65.000 246.820 ;
        END
    END VDDO
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        PORT
        LAYER M3 ;
        RECT  64.200 163.510 65.000 190.890 ;
        RECT  0.000 163.510 0.800 190.890 ;
        LAYER M2 ;
        RECT  0.000 172.080 65.000 183.060 ;
        LAYER TOP_M ;
        RECT  0.000 163.500 65.000 194.560 ;
        END
    END VDD
    PIN VSSO
        DIRECTION INOUT ;
        USE ground ;
        PORT
        LAYER M3 ;
        RECT  0.000 92.060 65.000 123.250 ;
        RECT  64.200 149.940 65.000 162.610 ;
        RECT  0.000 149.940 0.800 162.610 ;
        LAYER M2 ;
        RECT  0.000 147.040 65.000 154.520 ;
        LAYER TOP_M ;
        RECT  0.000 92.060 65.000 123.250 ;
        RECT  0.000 155.410 65.000 162.610 ;
        END
    END VSSO
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        PORT
        LAYER M3 ;
        RECT  64.200 130.690 65.000 148.880 ;
        RECT  0.000 130.690 0.800 148.880 ;
        LAYER M2 ;
        RECT  0.000 136.310 65.000 146.340 ;
        LAYER TOP_M ;
        RECT  0.000 123.850 65.000 154.560 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  2.000 0.000 63.000 250.000 ;
        RECT  0.000 88.990 65.000 130.360 ;
        RECT  0.000 136.510 65.000 157.550 ;
        RECT  0.315 158.150 64.700 158.460 ;
        RECT  0.300 158.930 64.700 159.230 ;
        RECT  0.300 159.530 64.700 159.830 ;
        RECT  0.300 160.130 64.700 160.430 ;
        RECT  0.300 160.730 64.700 161.030 ;
        RECT  0.300 161.330 64.700 161.630 ;
        RECT  0.300 161.910 64.700 162.190 ;
        RECT  0.300 162.490 64.700 162.770 ;
        RECT  0.300 163.070 64.700 163.350 ;
        RECT  0.300 163.650 64.700 163.950 ;
        RECT  0.300 164.250 64.700 164.550 ;
        RECT  0.300 164.850 64.700 165.150 ;
        RECT  0.300 165.450 64.700 165.750 ;
        RECT  0.300 166.050 64.700 166.350 ;
        RECT  0.300 166.650 64.700 166.960 ;
        RECT  0.300 167.260 64.700 167.560 ;
        RECT  0.300 167.860 64.700 168.160 ;
        RECT  0.000 169.150 65.000 197.240 ;
        RECT  0.600 0.600 64.400 250.000 ;
        RECT  0.000 198.470 65.000 250.000 ;
        LAYER M2 ;
        RECT  63.180 196.430 63.670 249.400 ;
        RECT  0.600 196.440 64.400 245.485 ;
        RECT  26.530 196.440 64.400 248.790 ;
        RECT  0.600 196.440 22.950 249.400 ;
        RECT  26.530 196.440 27.050 249.400 ;
        RECT  30.390 196.440 64.400 249.400 ;
        RECT  0.600 183.850 64.400 185.680 ;
        RECT  46.230 183.850 51.730 185.870 ;
        RECT  4.480 154.920 7.530 171.290 ;
        RECT  8.170 155.125 8.490 171.290 ;
        RECT  21.210 155.160 21.560 171.290 ;
        RECT  21.860 155.140 22.180 171.290 ;
        RECT  31.895 155.120 35.765 171.290 ;
        RECT  53.655 155.035 53.935 171.290 ;
        RECT  56.365 155.280 56.645 171.290 ;
        RECT  57.120 155.300 57.400 171.290 ;
        RECT  57.835 155.130 58.115 171.290 ;
        RECT  0.600 155.310 64.400 171.290 ;
        RECT  53.895 155.310 55.870 171.370 ;
        RECT  3.170 155.310 3.450 171.380 ;
        RECT  34.655 155.310 38.715 171.480 ;
        RECT  39.605 155.310 42.020 171.480 ;
        RECT  2.000 0.000 63.000 60.210 ;
        RECT  0.600 0.600 64.400 60.210 ;
        RECT  0.600 0.600 1.210 135.520 ;
        RECT  0.600 91.020 64.400 135.520 ;
        RECT  4.080 91.020 60.940 135.690 ;
        RECT  62.580 91.020 62.995 135.710 ;
        LAYER M3 ;
        RECT  0.600 247.660 23.220 248.740 ;
        RECT  0.600 247.660 22.900 249.400 ;
        RECT  26.260 247.660 64.400 248.740 ;
        RECT  26.580 247.660 27.000 249.400 ;
        RECT  30.440 247.660 64.400 249.400 ;
        RECT  0.600 124.090 64.400 129.850 ;
        RECT  1.640 124.090 63.600 135.790 ;
        RECT  1.810 124.090 2.830 154.520 ;
        RECT  3.510 124.090 63.600 171.560 ;
        RECT  4.040 123.970 60.900 171.560 ;
        RECT  1.640 155.040 63.600 171.560 ;
        RECT  1.640 183.580 63.600 185.950 ;
        RECT  5.515 124.090 63.600 200.820 ;
        RECT  1.640 196.170 63.600 200.820 ;
        RECT  0.600 0.600 64.400 60.480 ;
        RECT  2.000 0.000 63.000 88.700 ;
        RECT  0.600 0.600 1.480 91.220 ;
        RECT  0.600 90.750 64.400 91.220 ;
        LAYER TOP_M ;
        RECT  0.600 247.690 64.400 248.850 ;
        RECT  0.600 247.690 23.010 249.400 ;
        RECT  26.470 247.690 27.110 249.400 ;
        RECT  30.330 247.690 64.400 249.400 ;
        RECT  2.000 0.000 63.000 91.190 ;
        RECT  0.600 0.600 64.400 91.190 ;
    END
END pt3t03

MACRO pt3t02u
    CLASS PAD ;
    FOREIGN pt3t02u 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 65.000 BY 250.000 ;
    SYMMETRY X Y R90 ;
    SITE IOSite_c ;
    PIN PAD
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 55.440  LAYER TOP_M  ;
        ANTENNAPARTIALMETALSIDEAREA 287.938  LAYER M3  ;
        ANTENNAPARTIALMETALSIDEAREA 480.740  LAYER M2  ;
        ANTENNADIFFAREA 2657.280  LAYER TOP_M  ;
        ANTENNADIFFAREA 2657.280  LAYER M3  ;
        ANTENNADIFFAREA 1209.600  LAYER M2  ;
        ANTENNAPARTIALCUTAREA 632.318  LAYER TOP_V  ;
        ANTENNAPARTIALCUTAREA 349.898  LAYER V3  ;
        ANTENNAPARTIALCUTAREA 255.798  LAYER V2  ;
        PORT
        LAYER M3 ;
        RECT  23.740 249.580 25.740 250.000 ;
        LAYER M2 ;
        RECT  2.000 61.000 63.000 90.230 ;
        RECT  23.740 246.275 25.740 250.000 ;
        END
    END PAD
    PIN OEN
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 67.374  LAYER M1  ;
        ANTENNAPARTIALMETALSIDEAREA 81.726  LAYER M2  ;
        ANTENNAPARTIALMETALSIDEAREA 41.679  LAYER M3  ;
        ANTENNADIFFAREA 0.250  LAYER M3  ;
        ANTENNAPARTIALCUTAREA 0.203  LAYER V2  ;
        ANTENNAPARTIALCUTAREA 0.135  LAYER V3  ;
        ANTENNAGATEAREA 8.100  LAYER M2  ;
        ANTENNAGATEAREA 9.900  LAYER M3  ;
        PORT
        LAYER M3 ;
        RECT  28.870 249.580 29.600 250.000 ;
        LAYER M2 ;
        RECT  28.870 249.580 29.600 250.000 ;
        END
    END OEN
    PIN I
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 80.804  LAYER M2  ;
        ANTENNAPARTIALMETALSIDEAREA 67.374  LAYER M1  ;
        ANTENNAPARTIALMETALSIDEAREA 41.096  LAYER M3  ;
        ANTENNADIFFAREA 0.250  LAYER M3  ;
        ANTENNAPARTIALCUTAREA 0.135  LAYER V3  ;
        ANTENNAPARTIALCUTAREA 0.270  LAYER V2  ;
        ANTENNAGATEAREA 18.900  LAYER M2  ;
        ANTENNAGATEAREA 20.700  LAYER M3  ;
        PORT
        LAYER M3 ;
        RECT  27.840 249.580 28.570 250.000 ;
        LAYER M2 ;
        RECT  27.840 249.580 28.570 250.000 ;
        END
    END I
    PIN VDDO
        DIRECTION INOUT ;
        USE power ;
        PORT
        LAYER M3 ;
        RECT  64.200 192.330 65.000 200.640 ;
        RECT  0.000 201.660 65.000 221.520 ;
        RECT  0.000 222.720 65.000 246.820 ;
        RECT  0.000 192.330 0.800 200.640 ;
        LAYER M2 ;
        RECT  0.000 186.470 65.000 195.650 ;
        LAYER TOP_M ;
        RECT  0.000 195.170 65.000 200.640 ;
        RECT  0.000 201.660 65.000 221.520 ;
        RECT  0.000 222.720 65.000 246.820 ;
        END
    END VDDO
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        PORT
        LAYER M3 ;
        RECT  64.200 163.510 65.000 190.890 ;
        RECT  0.000 163.510 0.800 190.890 ;
        LAYER M2 ;
        RECT  0.000 172.080 65.000 183.060 ;
        LAYER TOP_M ;
        RECT  0.000 163.500 65.000 194.560 ;
        END
    END VDD
    PIN VSSO
        DIRECTION INOUT ;
        USE ground ;
        PORT
        LAYER M3 ;
        RECT  0.000 92.060 65.000 123.250 ;
        RECT  64.200 149.940 65.000 162.610 ;
        RECT  0.000 149.940 0.800 162.610 ;
        LAYER M2 ;
        RECT  0.000 147.040 65.000 154.520 ;
        LAYER TOP_M ;
        RECT  0.000 92.060 65.000 123.250 ;
        RECT  0.000 155.410 65.000 162.610 ;
        END
    END VSSO
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        PORT
        LAYER M3 ;
        RECT  64.200 130.690 65.000 148.880 ;
        RECT  0.000 130.690 0.800 148.880 ;
        LAYER M2 ;
        RECT  0.000 136.310 65.000 146.340 ;
        LAYER TOP_M ;
        RECT  0.000 123.850 65.000 154.560 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  2.000 0.000 63.000 250.000 ;
        RECT  0.000 88.990 65.000 130.360 ;
        RECT  0.000 136.510 65.000 157.550 ;
        RECT  0.315 158.150 64.700 158.460 ;
        RECT  0.300 158.930 64.700 159.230 ;
        RECT  0.300 159.530 64.700 159.830 ;
        RECT  0.300 160.130 64.700 160.430 ;
        RECT  0.300 160.730 64.700 161.030 ;
        RECT  0.300 161.330 64.700 161.630 ;
        RECT  0.300 161.910 64.700 162.190 ;
        RECT  0.300 162.490 64.700 162.770 ;
        RECT  0.300 163.070 64.700 163.350 ;
        RECT  0.300 163.650 64.700 163.950 ;
        RECT  0.300 164.250 64.700 164.550 ;
        RECT  0.300 164.850 64.700 165.150 ;
        RECT  0.300 165.450 64.700 165.750 ;
        RECT  0.300 166.050 64.700 166.350 ;
        RECT  0.300 166.650 64.700 166.960 ;
        RECT  0.300 167.260 64.700 167.560 ;
        RECT  0.300 167.860 64.700 168.160 ;
        RECT  0.000 169.150 65.000 197.240 ;
        RECT  0.600 0.600 64.400 250.000 ;
        RECT  0.000 198.470 65.000 250.000 ;
        LAYER M2 ;
        RECT  63.180 196.430 63.670 249.400 ;
        RECT  0.600 196.440 64.400 245.485 ;
        RECT  26.530 196.440 64.400 248.790 ;
        RECT  0.600 196.440 22.950 249.400 ;
        RECT  26.530 196.440 27.050 249.400 ;
        RECT  30.390 196.440 64.400 249.400 ;
        RECT  0.600 183.850 64.400 185.680 ;
        RECT  46.230 183.850 51.730 185.870 ;
        RECT  4.895 155.120 7.525 171.290 ;
        RECT  8.170 155.125 8.490 171.290 ;
        RECT  21.080 155.160 21.430 171.290 ;
        RECT  21.730 155.140 22.050 171.290 ;
        RECT  53.655 155.035 53.935 171.290 ;
        RECT  56.365 155.280 56.645 171.290 ;
        RECT  57.120 155.300 57.400 171.290 ;
        RECT  57.835 155.130 58.115 171.290 ;
        RECT  0.600 155.310 64.400 171.290 ;
        RECT  53.895 155.310 55.870 171.370 ;
        RECT  33.190 155.310 33.690 171.375 ;
        RECT  3.210 155.310 3.490 171.380 ;
        RECT  34.655 155.310 38.715 171.480 ;
        RECT  39.605 155.310 42.020 171.480 ;
        RECT  2.000 0.000 63.000 60.210 ;
        RECT  0.600 0.600 64.400 60.210 ;
        RECT  0.600 0.600 1.210 135.520 ;
        RECT  0.600 91.020 64.400 135.520 ;
        RECT  4.080 91.020 60.940 135.690 ;
        RECT  62.580 91.020 62.995 135.710 ;
        LAYER M3 ;
        RECT  0.600 247.660 23.220 248.740 ;
        RECT  0.600 247.660 22.900 249.400 ;
        RECT  26.260 247.660 64.400 248.740 ;
        RECT  26.580 247.660 27.000 249.400 ;
        RECT  30.440 247.660 64.400 249.400 ;
        RECT  0.600 124.090 64.400 129.850 ;
        RECT  1.640 124.090 63.600 135.790 ;
        RECT  1.810 124.090 2.830 154.520 ;
        RECT  3.110 124.090 63.600 171.560 ;
        RECT  4.040 123.970 60.900 171.560 ;
        RECT  1.640 155.040 63.600 171.560 ;
        RECT  1.640 183.580 63.600 185.950 ;
        RECT  5.510 124.090 63.600 200.820 ;
        RECT  1.640 196.170 63.600 200.820 ;
        RECT  0.600 0.600 64.400 60.480 ;
        RECT  2.000 0.000 63.000 88.700 ;
        RECT  0.600 0.600 1.480 91.220 ;
        RECT  0.600 90.750 64.400 91.220 ;
        LAYER TOP_M ;
        RECT  0.600 247.690 64.400 248.850 ;
        RECT  0.600 247.690 23.010 249.400 ;
        RECT  26.470 247.690 27.110 249.400 ;
        RECT  30.330 247.690 64.400 249.400 ;
        RECT  2.000 0.000 63.000 91.190 ;
        RECT  0.600 0.600 64.400 91.190 ;
    END
END pt3t02u

MACRO pt3t02d
    CLASS PAD ;
    FOREIGN pt3t02d 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 65.000 BY 250.000 ;
    SYMMETRY X Y R90 ;
    SITE IOSite_c ;
    PIN PAD
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 55.440  LAYER TOP_M  ;
        ANTENNAPARTIALMETALSIDEAREA 287.938  LAYER M3  ;
        ANTENNAPARTIALMETALSIDEAREA 480.740  LAYER M2  ;
        ANTENNADIFFAREA 2657.280  LAYER TOP_M  ;
        ANTENNADIFFAREA 2657.280  LAYER M3  ;
        ANTENNADIFFAREA 1209.600  LAYER M2  ;
        ANTENNAPARTIALCUTAREA 632.318  LAYER TOP_V  ;
        ANTENNAPARTIALCUTAREA 349.898  LAYER V3  ;
        ANTENNAPARTIALCUTAREA 255.798  LAYER V2  ;
        PORT
        LAYER M3 ;
        RECT  23.740 249.580 25.740 250.000 ;
        LAYER M2 ;
        RECT  2.000 61.000 63.000 90.230 ;
        RECT  23.740 246.275 25.740 250.000 ;
        END
    END PAD
    PIN OEN
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 81.726  LAYER M2  ;
        ANTENNAPARTIALMETALSIDEAREA 67.374  LAYER M1  ;
        ANTENNAPARTIALMETALSIDEAREA 41.679  LAYER M3  ;
        ANTENNADIFFAREA 0.250  LAYER M3  ;
        ANTENNAPARTIALCUTAREA 0.203  LAYER V2  ;
        ANTENNAPARTIALCUTAREA 0.135  LAYER V3  ;
        ANTENNAGATEAREA 8.100  LAYER M2  ;
        ANTENNAGATEAREA 9.900  LAYER M3  ;
        PORT
        LAYER M3 ;
        RECT  28.870 249.580 29.600 250.000 ;
        LAYER M2 ;
        RECT  28.870 249.580 29.600 250.000 ;
        END
    END OEN
    PIN I
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 67.374  LAYER M1  ;
        ANTENNAPARTIALMETALSIDEAREA 80.804  LAYER M2  ;
        ANTENNAPARTIALMETALSIDEAREA 41.096  LAYER M3  ;
        ANTENNADIFFAREA 0.250  LAYER M3  ;
        ANTENNAPARTIALCUTAREA 0.270  LAYER V2  ;
        ANTENNAPARTIALCUTAREA 0.135  LAYER V3  ;
        ANTENNAGATEAREA 18.900  LAYER M2  ;
        ANTENNAGATEAREA 20.700  LAYER M3  ;
        PORT
        LAYER M3 ;
        RECT  27.840 249.580 28.570 250.000 ;
        LAYER M2 ;
        RECT  27.840 249.580 28.570 250.000 ;
        END
    END I
    PIN VDDO
        DIRECTION INOUT ;
        USE power ;
        PORT
        LAYER M3 ;
        RECT  64.200 192.330 65.000 200.640 ;
        RECT  0.000 201.660 65.000 221.520 ;
        RECT  0.000 222.720 65.000 246.820 ;
        RECT  0.000 192.330 0.800 200.640 ;
        LAYER M2 ;
        RECT  0.000 186.470 65.000 195.650 ;
        LAYER TOP_M ;
        RECT  0.000 195.170 65.000 200.640 ;
        RECT  0.000 201.660 65.000 221.520 ;
        RECT  0.000 222.720 65.000 246.820 ;
        END
    END VDDO
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        PORT
        LAYER M3 ;
        RECT  64.200 163.510 65.000 190.890 ;
        RECT  0.000 163.510 0.800 190.890 ;
        LAYER M2 ;
        RECT  0.000 172.080 65.000 183.060 ;
        LAYER TOP_M ;
        RECT  0.000 163.500 65.000 194.560 ;
        END
    END VDD
    PIN VSSO
        DIRECTION INOUT ;
        USE ground ;
        PORT
        LAYER M3 ;
        RECT  0.000 92.060 65.000 123.250 ;
        RECT  64.200 149.940 65.000 162.610 ;
        RECT  0.000 149.940 0.800 162.610 ;
        LAYER M2 ;
        RECT  0.000 147.040 65.000 154.520 ;
        LAYER TOP_M ;
        RECT  0.000 92.060 65.000 123.250 ;
        RECT  0.000 155.410 65.000 162.610 ;
        END
    END VSSO
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        PORT
        LAYER M3 ;
        RECT  64.200 130.690 65.000 148.880 ;
        RECT  0.000 130.690 0.800 148.880 ;
        LAYER M2 ;
        RECT  0.000 136.310 65.000 146.340 ;
        LAYER TOP_M ;
        RECT  0.000 123.850 65.000 154.560 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  2.000 0.000 63.000 250.000 ;
        RECT  0.000 88.990 65.000 130.360 ;
        RECT  0.000 136.510 65.000 157.550 ;
        RECT  0.315 158.150 64.700 158.460 ;
        RECT  0.300 158.930 64.700 159.230 ;
        RECT  0.300 159.530 64.700 159.830 ;
        RECT  0.300 160.130 64.700 160.430 ;
        RECT  0.300 160.730 64.700 161.030 ;
        RECT  0.300 161.330 64.700 161.630 ;
        RECT  0.300 161.910 64.700 162.190 ;
        RECT  0.300 162.490 64.700 162.770 ;
        RECT  0.300 163.070 64.700 163.350 ;
        RECT  0.300 163.650 64.700 163.950 ;
        RECT  0.300 164.250 64.700 164.550 ;
        RECT  0.300 164.850 64.700 165.150 ;
        RECT  0.300 165.450 64.700 165.750 ;
        RECT  0.300 166.050 64.700 166.350 ;
        RECT  0.300 166.650 64.700 166.960 ;
        RECT  0.300 167.260 64.700 167.560 ;
        RECT  0.300 167.860 64.700 168.160 ;
        RECT  0.000 169.150 65.000 197.240 ;
        RECT  0.600 0.600 64.400 250.000 ;
        RECT  0.000 198.470 65.000 250.000 ;
        LAYER M2 ;
        RECT  63.180 196.430 63.670 249.400 ;
        RECT  0.600 196.440 64.400 245.485 ;
        RECT  26.530 196.440 64.400 248.790 ;
        RECT  0.600 196.440 22.950 249.400 ;
        RECT  26.530 196.440 27.050 249.400 ;
        RECT  30.390 196.440 64.400 249.400 ;
        RECT  0.600 183.850 64.400 185.680 ;
        RECT  46.230 183.850 51.730 185.870 ;
        RECT  4.895 155.120 7.525 171.290 ;
        RECT  8.170 155.125 8.490 171.290 ;
        RECT  21.080 155.160 21.430 171.290 ;
        RECT  21.730 155.140 22.050 171.290 ;
        RECT  49.115 155.130 51.355 171.290 ;
        RECT  52.295 155.300 52.605 171.290 ;
        RECT  53.655 155.035 53.935 171.290 ;
        RECT  56.365 155.280 56.645 171.290 ;
        RECT  57.120 155.300 57.400 171.290 ;
        RECT  57.835 155.130 58.115 171.290 ;
        RECT  0.600 155.310 64.400 171.290 ;
        RECT  53.895 155.310 55.870 171.370 ;
        RECT  3.210 155.310 3.490 171.380 ;
        RECT  34.655 155.310 38.715 171.480 ;
        RECT  39.605 155.310 42.020 171.480 ;
        RECT  2.000 0.000 63.000 60.210 ;
        RECT  0.600 0.600 64.400 60.210 ;
        RECT  0.600 0.600 1.210 135.520 ;
        RECT  0.600 91.020 64.400 135.520 ;
        RECT  4.080 91.020 60.940 135.690 ;
        RECT  62.580 91.020 62.995 135.710 ;
        LAYER M3 ;
        RECT  0.600 247.660 23.220 248.740 ;
        RECT  0.600 247.660 22.900 249.400 ;
        RECT  26.260 247.660 64.400 248.740 ;
        RECT  26.580 247.660 27.000 249.400 ;
        RECT  30.440 247.660 64.400 249.400 ;
        RECT  0.600 124.090 64.400 129.850 ;
        RECT  1.640 124.090 63.600 135.790 ;
        RECT  1.810 124.090 2.830 154.520 ;
        RECT  3.110 124.090 63.600 171.560 ;
        RECT  4.040 123.970 60.900 171.560 ;
        RECT  1.640 155.040 63.600 171.560 ;
        RECT  1.640 183.580 63.600 185.950 ;
        RECT  5.510 124.090 63.600 200.820 ;
        RECT  1.640 196.170 63.600 200.820 ;
        RECT  0.600 0.600 64.400 60.480 ;
        RECT  2.000 0.000 63.000 88.700 ;
        RECT  0.600 0.600 1.480 91.220 ;
        RECT  0.600 90.750 64.400 91.220 ;
        LAYER TOP_M ;
        RECT  0.600 247.690 64.400 248.850 ;
        RECT  0.600 247.690 23.010 249.400 ;
        RECT  26.470 247.690 27.110 249.400 ;
        RECT  30.330 247.690 64.400 249.400 ;
        RECT  2.000 0.000 63.000 91.190 ;
        RECT  0.600 0.600 64.400 91.190 ;
    END
END pt3t02d

MACRO pt3t02
    CLASS PAD ;
    FOREIGN pt3t02 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 65.000 BY 250.000 ;
    SYMMETRY X Y R90 ;
    SITE IOSite_c ;
    PIN PAD
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 55.440  LAYER TOP_M  ;
        ANTENNAPARTIALMETALSIDEAREA 287.938  LAYER M3  ;
        ANTENNAPARTIALMETALSIDEAREA 480.740  LAYER M2  ;
        ANTENNADIFFAREA 2657.280  LAYER TOP_M  ;
        ANTENNADIFFAREA 2657.280  LAYER M3  ;
        ANTENNADIFFAREA 1209.600  LAYER M2  ;
        ANTENNAPARTIALCUTAREA 632.318  LAYER TOP_V  ;
        ANTENNAPARTIALCUTAREA 349.898  LAYER V3  ;
        ANTENNAPARTIALCUTAREA 255.798  LAYER V2  ;
        PORT
        LAYER M3 ;
        RECT  23.740 249.580 25.740 250.000 ;
        LAYER M2 ;
        RECT  2.000 61.000 63.000 90.230 ;
        RECT  23.740 246.275 25.740 250.000 ;
        END
    END PAD
    PIN OEN
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 67.374  LAYER M1  ;
        ANTENNAPARTIALMETALSIDEAREA 81.726  LAYER M2  ;
        ANTENNAPARTIALMETALSIDEAREA 41.679  LAYER M3  ;
        ANTENNADIFFAREA 0.250  LAYER M3  ;
        ANTENNAPARTIALCUTAREA 0.203  LAYER V2  ;
        ANTENNAPARTIALCUTAREA 0.135  LAYER V3  ;
        ANTENNAGATEAREA 8.100  LAYER M2  ;
        ANTENNAGATEAREA 9.900  LAYER M3  ;
        PORT
        LAYER M3 ;
        RECT  28.870 249.580 29.600 250.000 ;
        LAYER M2 ;
        RECT  28.870 249.580 29.600 250.000 ;
        END
    END OEN
    PIN I
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 67.374  LAYER M1  ;
        ANTENNAPARTIALMETALSIDEAREA 80.804  LAYER M2  ;
        ANTENNAPARTIALMETALSIDEAREA 41.096  LAYER M3  ;
        ANTENNADIFFAREA 0.250  LAYER M3  ;
        ANTENNAPARTIALCUTAREA 0.270  LAYER V2  ;
        ANTENNAPARTIALCUTAREA 0.135  LAYER V3  ;
        ANTENNAGATEAREA 18.900  LAYER M2  ;
        ANTENNAGATEAREA 20.700  LAYER M3  ;
        PORT
        LAYER M3 ;
        RECT  27.840 249.580 28.570 250.000 ;
        LAYER M2 ;
        RECT  27.840 249.580 28.570 250.000 ;
        END
    END I
    PIN VDDO
        DIRECTION INOUT ;
        USE power ;
        PORT
        LAYER M3 ;
        RECT  64.200 192.330 65.000 200.640 ;
        RECT  0.000 201.660 65.000 221.520 ;
        RECT  0.000 222.720 65.000 246.820 ;
        RECT  0.000 192.330 0.800 200.640 ;
        LAYER M2 ;
        RECT  0.000 186.470 65.000 195.650 ;
        LAYER TOP_M ;
        RECT  0.000 195.170 65.000 200.640 ;
        RECT  0.000 201.660 65.000 221.520 ;
        RECT  0.000 222.720 65.000 246.820 ;
        END
    END VDDO
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        PORT
        LAYER M3 ;
        RECT  64.200 163.510 65.000 190.890 ;
        RECT  0.000 163.510 0.800 190.890 ;
        LAYER M2 ;
        RECT  0.000 172.080 65.000 183.060 ;
        LAYER TOP_M ;
        RECT  0.000 163.500 65.000 194.560 ;
        END
    END VDD
    PIN VSSO
        DIRECTION INOUT ;
        USE ground ;
        PORT
        LAYER M3 ;
        RECT  0.000 92.060 65.000 123.250 ;
        RECT  64.200 149.940 65.000 162.610 ;
        RECT  0.000 149.940 0.800 162.610 ;
        LAYER M2 ;
        RECT  0.000 147.040 65.000 154.520 ;
        LAYER TOP_M ;
        RECT  0.000 92.060 65.000 123.250 ;
        RECT  0.000 155.410 65.000 162.610 ;
        END
    END VSSO
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        PORT
        LAYER M3 ;
        RECT  64.200 130.690 65.000 148.880 ;
        RECT  0.000 130.690 0.800 148.880 ;
        LAYER M2 ;
        RECT  0.000 136.310 65.000 146.340 ;
        LAYER TOP_M ;
        RECT  0.000 123.850 65.000 154.560 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  2.000 0.000 63.000 250.000 ;
        RECT  0.000 88.990 65.000 130.360 ;
        RECT  0.000 136.510 65.000 157.550 ;
        RECT  0.315 158.150 64.700 158.460 ;
        RECT  0.300 158.930 64.700 159.230 ;
        RECT  0.300 159.530 64.700 159.830 ;
        RECT  0.300 160.130 64.700 160.430 ;
        RECT  0.300 160.730 64.700 161.030 ;
        RECT  0.300 161.330 64.700 161.630 ;
        RECT  0.300 161.910 64.700 162.190 ;
        RECT  0.300 162.490 64.700 162.770 ;
        RECT  0.300 163.070 64.700 163.350 ;
        RECT  0.300 163.650 64.700 163.950 ;
        RECT  0.300 164.250 64.700 164.550 ;
        RECT  0.300 164.850 64.700 165.150 ;
        RECT  0.300 165.450 64.700 165.750 ;
        RECT  0.300 166.050 64.700 166.350 ;
        RECT  0.300 166.650 64.700 166.960 ;
        RECT  0.300 167.260 64.700 167.560 ;
        RECT  0.300 167.860 64.700 168.160 ;
        RECT  0.000 169.150 65.000 197.240 ;
        RECT  0.600 0.600 64.400 250.000 ;
        RECT  0.000 198.470 65.000 250.000 ;
        LAYER M2 ;
        RECT  63.180 196.430 63.670 249.400 ;
        RECT  0.600 196.440 64.400 245.485 ;
        RECT  26.530 196.440 64.400 248.790 ;
        RECT  0.600 196.440 22.950 249.400 ;
        RECT  26.530 196.440 27.050 249.400 ;
        RECT  30.390 196.440 64.400 249.400 ;
        RECT  0.600 183.850 64.400 185.680 ;
        RECT  46.230 183.850 51.730 185.870 ;
        RECT  4.895 155.120 7.525 171.290 ;
        RECT  8.170 155.125 8.490 171.290 ;
        RECT  21.080 155.160 21.430 171.290 ;
        RECT  21.730 155.140 22.050 171.290 ;
        RECT  53.655 155.035 53.935 171.290 ;
        RECT  56.365 155.280 56.645 171.290 ;
        RECT  57.120 155.300 57.400 171.290 ;
        RECT  57.835 155.130 58.115 171.290 ;
        RECT  0.600 155.310 64.400 171.290 ;
        RECT  53.895 155.310 55.870 171.370 ;
        RECT  3.210 155.310 3.490 171.380 ;
        RECT  34.655 155.310 38.715 171.480 ;
        RECT  39.605 155.310 42.020 171.480 ;
        RECT  2.000 0.000 63.000 60.210 ;
        RECT  0.600 0.600 64.400 60.210 ;
        RECT  0.600 0.600 1.210 135.520 ;
        RECT  0.600 91.020 64.400 135.520 ;
        RECT  4.080 91.020 60.940 135.690 ;
        RECT  62.580 91.020 62.995 135.710 ;
        LAYER M3 ;
        RECT  0.600 247.660 23.220 248.740 ;
        RECT  0.600 247.660 22.900 249.400 ;
        RECT  26.260 247.660 64.400 248.740 ;
        RECT  26.580 247.660 27.000 249.400 ;
        RECT  30.440 247.660 64.400 249.400 ;
        RECT  0.600 124.090 64.400 129.850 ;
        RECT  1.640 124.090 63.600 135.790 ;
        RECT  1.810 124.090 2.830 154.520 ;
        RECT  3.110 124.090 63.600 171.560 ;
        RECT  4.040 123.970 60.900 171.560 ;
        RECT  1.640 155.040 63.600 171.560 ;
        RECT  1.640 183.580 63.600 185.950 ;
        RECT  5.510 124.090 63.600 200.820 ;
        RECT  1.640 196.170 63.600 200.820 ;
        RECT  0.600 0.600 64.400 60.480 ;
        RECT  2.000 0.000 63.000 88.700 ;
        RECT  0.600 0.600 1.480 91.220 ;
        RECT  0.600 90.750 64.400 91.220 ;
        LAYER TOP_M ;
        RECT  0.600 247.690 64.400 248.850 ;
        RECT  0.600 247.690 23.010 249.400 ;
        RECT  26.470 247.690 27.110 249.400 ;
        RECT  30.330 247.690 64.400 249.400 ;
        RECT  2.000 0.000 63.000 91.190 ;
        RECT  0.600 0.600 64.400 91.190 ;
    END
END pt3t02

MACRO pt3t01u
    CLASS PAD ;
    FOREIGN pt3t01u 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 65.000 BY 250.000 ;
    SYMMETRY X Y R90 ;
    SITE IOSite_c ;
    PIN PAD
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 55.440  LAYER TOP_M  ;
        ANTENNAPARTIALMETALSIDEAREA 287.938  LAYER M3  ;
        ANTENNAPARTIALMETALSIDEAREA 480.740  LAYER M2  ;
        ANTENNADIFFAREA 2657.280  LAYER TOP_M  ;
        ANTENNADIFFAREA 2657.280  LAYER M3  ;
        ANTENNADIFFAREA 1209.600  LAYER M2  ;
        ANTENNAPARTIALCUTAREA 632.318  LAYER TOP_V  ;
        ANTENNAPARTIALCUTAREA 349.898  LAYER V3  ;
        ANTENNAPARTIALCUTAREA 255.798  LAYER V2  ;
        PORT
        LAYER M3 ;
        RECT  23.740 249.580 25.740 250.000 ;
        LAYER M2 ;
        RECT  2.000 61.000 63.000 90.230 ;
        RECT  23.740 246.275 25.740 250.000 ;
        END
    END PAD
    PIN OEN
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 81.726  LAYER M2  ;
        ANTENNAPARTIALMETALSIDEAREA 67.374  LAYER M1  ;
        ANTENNAPARTIALMETALSIDEAREA 41.679  LAYER M3  ;
        ANTENNADIFFAREA 0.250  LAYER M3  ;
        ANTENNAPARTIALCUTAREA 0.203  LAYER V2  ;
        ANTENNAPARTIALCUTAREA 0.135  LAYER V3  ;
        ANTENNAGATEAREA 8.100  LAYER M2  ;
        ANTENNAGATEAREA 9.900  LAYER M3  ;
        PORT
        LAYER M3 ;
        RECT  28.870 249.580 29.600 250.000 ;
        LAYER M2 ;
        RECT  28.870 249.580 29.600 250.000 ;
        END
    END OEN
    PIN I
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 67.374  LAYER M1  ;
        ANTENNAPARTIALMETALSIDEAREA 80.804  LAYER M2  ;
        ANTENNAPARTIALMETALSIDEAREA 41.096  LAYER M3  ;
        ANTENNADIFFAREA 0.250  LAYER M3  ;
        ANTENNAPARTIALCUTAREA 0.203  LAYER V2  ;
        ANTENNAPARTIALCUTAREA 0.135  LAYER V3  ;
        ANTENNAGATEAREA 8.100  LAYER M2  ;
        ANTENNAGATEAREA 9.900  LAYER M3  ;
        PORT
        LAYER M3 ;
        RECT  27.840 249.580 28.570 250.000 ;
        LAYER M2 ;
        RECT  27.840 249.580 28.570 250.000 ;
        END
    END I
    PIN VDDO
        DIRECTION INOUT ;
        USE power ;
        PORT
        LAYER M3 ;
        RECT  64.200 192.330 65.000 200.640 ;
        RECT  0.000 201.660 65.000 221.520 ;
        RECT  0.000 222.720 65.000 246.820 ;
        RECT  0.000 192.330 0.800 200.640 ;
        LAYER M2 ;
        RECT  0.000 186.470 65.000 195.650 ;
        LAYER TOP_M ;
        RECT  0.000 195.170 65.000 200.640 ;
        RECT  0.000 201.660 65.000 221.520 ;
        RECT  0.000 222.720 65.000 246.820 ;
        END
    END VDDO
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        PORT
        LAYER M3 ;
        RECT  64.200 163.510 65.000 190.890 ;
        RECT  0.000 163.510 0.800 190.890 ;
        LAYER M2 ;
        RECT  0.000 172.080 65.000 183.060 ;
        LAYER TOP_M ;
        RECT  0.000 163.500 65.000 194.560 ;
        END
    END VDD
    PIN VSSO
        DIRECTION INOUT ;
        USE ground ;
        PORT
        LAYER M3 ;
        RECT  0.000 92.060 65.000 123.250 ;
        RECT  64.200 149.940 65.000 162.610 ;
        RECT  0.000 149.940 0.800 162.610 ;
        LAYER M2 ;
        RECT  0.000 147.040 65.000 154.520 ;
        LAYER TOP_M ;
        RECT  0.000 92.060 65.000 123.250 ;
        RECT  0.000 155.410 65.000 162.610 ;
        END
    END VSSO
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        PORT
        LAYER M3 ;
        RECT  64.200 130.690 65.000 148.880 ;
        RECT  0.000 130.690 0.800 148.880 ;
        LAYER M2 ;
        RECT  0.000 136.310 65.000 146.340 ;
        LAYER TOP_M ;
        RECT  0.000 123.850 65.000 154.560 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  2.000 0.000 63.000 250.000 ;
        RECT  0.000 88.990 65.000 130.360 ;
        RECT  0.000 136.510 65.000 157.550 ;
        RECT  0.315 158.150 64.700 158.460 ;
        RECT  0.300 158.930 64.700 159.230 ;
        RECT  0.300 159.530 64.700 159.830 ;
        RECT  0.300 160.130 64.700 160.430 ;
        RECT  0.300 160.730 64.700 161.030 ;
        RECT  0.300 161.330 64.700 161.630 ;
        RECT  0.300 161.910 64.700 162.190 ;
        RECT  0.300 162.490 64.700 162.770 ;
        RECT  0.300 163.070 64.700 163.350 ;
        RECT  0.300 163.650 64.700 163.950 ;
        RECT  0.300 164.250 64.700 164.550 ;
        RECT  0.300 164.850 64.700 165.150 ;
        RECT  0.300 165.450 64.700 165.750 ;
        RECT  0.300 166.050 64.700 166.350 ;
        RECT  0.300 166.650 64.700 166.960 ;
        RECT  0.300 167.260 64.700 167.560 ;
        RECT  0.300 167.860 64.700 168.160 ;
        RECT  0.000 169.150 65.000 197.240 ;
        RECT  0.600 0.600 64.400 250.000 ;
        RECT  0.000 198.470 65.000 250.000 ;
        LAYER M2 ;
        RECT  63.180 196.430 63.670 249.400 ;
        RECT  0.600 196.440 64.400 245.485 ;
        RECT  26.530 196.440 64.400 248.790 ;
        RECT  0.600 196.440 22.950 249.400 ;
        RECT  26.530 196.440 27.050 249.400 ;
        RECT  30.390 196.440 64.400 249.400 ;
        RECT  0.600 183.850 64.400 185.680 ;
        RECT  46.230 183.850 51.730 185.870 ;
        RECT  19.790 155.160 20.140 171.290 ;
        RECT  20.440 155.140 20.760 171.290 ;
        RECT  53.655 155.035 53.935 171.290 ;
        RECT  56.365 155.280 56.645 171.290 ;
        RECT  57.120 155.300 57.400 171.290 ;
        RECT  57.835 155.130 58.115 171.290 ;
        RECT  0.600 155.310 64.400 171.290 ;
        RECT  53.895 155.310 55.870 171.370 ;
        RECT  31.780 155.310 32.280 171.375 ;
        RECT  3.210 155.310 3.490 171.380 ;
        RECT  34.655 155.310 38.715 171.480 ;
        RECT  39.605 155.310 42.020 171.480 ;
        RECT  2.000 0.000 63.000 60.210 ;
        RECT  0.600 0.600 64.400 60.210 ;
        RECT  0.600 0.600 1.210 135.520 ;
        RECT  0.600 91.020 64.400 135.520 ;
        RECT  4.080 91.020 60.940 135.690 ;
        RECT  62.580 91.020 62.995 135.710 ;
        LAYER M3 ;
        RECT  0.600 247.660 23.220 248.740 ;
        RECT  0.600 247.660 22.900 249.400 ;
        RECT  26.260 247.660 64.400 248.740 ;
        RECT  26.580 247.660 27.000 249.400 ;
        RECT  30.440 247.660 64.400 249.400 ;
        RECT  0.600 124.090 64.400 129.850 ;
        RECT  3.990 123.970 60.900 135.790 ;
        RECT  1.640 124.090 63.600 135.790 ;
        RECT  1.810 124.090 2.830 154.520 ;
        RECT  5.155 123.970 60.900 171.560 ;
        RECT  1.640 155.040 63.600 171.560 ;
        RECT  1.640 183.580 63.600 185.950 ;
        RECT  5.490 124.090 63.600 200.820 ;
        RECT  1.640 196.170 63.600 200.820 ;
        RECT  0.600 0.600 64.400 60.480 ;
        RECT  2.000 0.000 63.000 88.700 ;
        RECT  0.600 0.600 1.480 91.220 ;
        RECT  0.600 90.750 64.400 91.220 ;
        LAYER TOP_M ;
        RECT  0.600 247.690 64.400 248.850 ;
        RECT  0.600 247.690 23.010 249.400 ;
        RECT  26.470 247.690 27.110 249.400 ;
        RECT  30.330 247.690 64.400 249.400 ;
        RECT  2.000 0.000 63.000 91.190 ;
        RECT  0.600 0.600 64.400 91.190 ;
    END
END pt3t01u

MACRO pt3t01d
    CLASS PAD ;
    FOREIGN pt3t01d 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 65.000 BY 250.000 ;
    SYMMETRY X Y R90 ;
    SITE IOSite_c ;
    PIN PAD
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 55.440  LAYER TOP_M  ;
        ANTENNAPARTIALMETALSIDEAREA 287.938  LAYER M3  ;
        ANTENNAPARTIALMETALSIDEAREA 480.740  LAYER M2  ;
        ANTENNADIFFAREA 2657.280  LAYER TOP_M  ;
        ANTENNADIFFAREA 2657.280  LAYER M3  ;
        ANTENNADIFFAREA 1209.600  LAYER M2  ;
        ANTENNAPARTIALCUTAREA 632.318  LAYER TOP_V  ;
        ANTENNAPARTIALCUTAREA 349.898  LAYER V3  ;
        ANTENNAPARTIALCUTAREA 255.798  LAYER V2  ;
        PORT
        LAYER M3 ;
        RECT  23.740 249.580 25.740 250.000 ;
        LAYER M2 ;
        RECT  2.000 61.000 63.000 90.230 ;
        RECT  23.740 246.275 25.740 250.000 ;
        END
    END PAD
    PIN OEN
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 81.726  LAYER M2  ;
        ANTENNAPARTIALMETALSIDEAREA 67.374  LAYER M1  ;
        ANTENNAPARTIALMETALSIDEAREA 41.679  LAYER M3  ;
        ANTENNADIFFAREA 0.250  LAYER M3  ;
        ANTENNAPARTIALCUTAREA 0.135  LAYER V3  ;
        ANTENNAPARTIALCUTAREA 0.203  LAYER V2  ;
        ANTENNAGATEAREA 8.100  LAYER M2  ;
        ANTENNAGATEAREA 9.900  LAYER M3  ;
        PORT
        LAYER M3 ;
        RECT  28.870 249.580 29.600 250.000 ;
        LAYER M2 ;
        RECT  28.870 249.580 29.600 250.000 ;
        END
    END OEN
    PIN I
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 80.804  LAYER M2  ;
        ANTENNAPARTIALMETALSIDEAREA 67.374  LAYER M1  ;
        ANTENNAPARTIALMETALSIDEAREA 41.096  LAYER M3  ;
        ANTENNADIFFAREA 0.250  LAYER M3  ;
        ANTENNAPARTIALCUTAREA 0.135  LAYER V3  ;
        ANTENNAPARTIALCUTAREA 0.203  LAYER V2  ;
        ANTENNAGATEAREA 8.100  LAYER M2  ;
        ANTENNAGATEAREA 9.900  LAYER M3  ;
        PORT
        LAYER M3 ;
        RECT  27.840 249.580 28.570 250.000 ;
        LAYER M2 ;
        RECT  27.840 249.580 28.570 250.000 ;
        END
    END I
    PIN VDDO
        DIRECTION INOUT ;
        USE power ;
        PORT
        LAYER M3 ;
        RECT  64.200 192.330 65.000 200.640 ;
        RECT  0.000 201.660 65.000 221.520 ;
        RECT  0.000 222.720 65.000 246.820 ;
        RECT  0.000 192.330 0.800 200.640 ;
        LAYER M2 ;
        RECT  0.000 186.470 65.000 195.650 ;
        LAYER TOP_M ;
        RECT  0.000 195.170 65.000 200.640 ;
        RECT  0.000 201.660 65.000 221.520 ;
        RECT  0.000 222.720 65.000 246.820 ;
        END
    END VDDO
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        PORT
        LAYER M3 ;
        RECT  64.200 163.510 65.000 190.890 ;
        RECT  0.000 163.510 0.800 190.890 ;
        LAYER M2 ;
        RECT  0.000 172.080 65.000 183.060 ;
        LAYER TOP_M ;
        RECT  0.000 163.500 65.000 194.560 ;
        END
    END VDD
    PIN VSSO
        DIRECTION INOUT ;
        USE ground ;
        PORT
        LAYER M3 ;
        RECT  0.000 92.060 65.000 123.250 ;
        RECT  64.200 149.940 65.000 162.610 ;
        RECT  0.000 149.940 0.800 162.610 ;
        LAYER M2 ;
        RECT  0.000 147.040 65.000 154.520 ;
        LAYER TOP_M ;
        RECT  0.000 92.060 65.000 123.250 ;
        RECT  0.000 155.410 65.000 162.610 ;
        END
    END VSSO
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        PORT
        LAYER M3 ;
        RECT  64.200 130.690 65.000 148.880 ;
        RECT  0.000 130.690 0.800 148.880 ;
        LAYER M2 ;
        RECT  0.000 136.310 65.000 146.340 ;
        LAYER TOP_M ;
        RECT  0.000 123.850 65.000 154.560 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  2.000 0.000 63.000 250.000 ;
        RECT  0.000 88.990 65.000 130.360 ;
        RECT  0.000 136.510 65.000 157.550 ;
        RECT  0.315 158.150 64.700 158.460 ;
        RECT  0.300 158.930 64.700 159.230 ;
        RECT  0.300 159.530 64.700 159.830 ;
        RECT  0.300 160.130 64.700 160.430 ;
        RECT  0.300 160.730 64.700 161.030 ;
        RECT  0.300 161.330 64.700 161.630 ;
        RECT  0.300 161.910 64.700 162.190 ;
        RECT  0.300 162.490 64.700 162.770 ;
        RECT  0.300 163.070 64.700 163.350 ;
        RECT  0.300 163.650 64.700 163.950 ;
        RECT  0.300 164.250 64.700 164.550 ;
        RECT  0.300 164.850 64.700 165.150 ;
        RECT  0.300 165.450 64.700 165.750 ;
        RECT  0.300 166.050 64.700 166.350 ;
        RECT  0.300 166.650 64.700 166.960 ;
        RECT  0.300 167.260 64.700 167.560 ;
        RECT  0.300 167.860 64.700 168.160 ;
        RECT  0.000 169.150 65.000 197.240 ;
        RECT  0.600 0.600 64.400 250.000 ;
        RECT  0.000 198.470 65.000 250.000 ;
        LAYER M2 ;
        RECT  63.180 196.430 63.670 249.400 ;
        RECT  0.600 196.440 64.400 245.485 ;
        RECT  26.530 196.440 64.400 248.790 ;
        RECT  0.600 196.440 22.950 249.400 ;
        RECT  26.530 196.440 27.050 249.400 ;
        RECT  30.390 196.440 64.400 249.400 ;
        RECT  0.600 183.850 64.400 185.680 ;
        RECT  46.230 183.850 51.730 185.870 ;
        RECT  19.790 155.160 20.140 171.290 ;
        RECT  20.440 155.140 20.760 171.290 ;
        RECT  49.330 155.130 51.570 171.290 ;
        RECT  52.510 155.300 52.820 171.290 ;
        RECT  53.655 155.035 53.935 171.290 ;
        RECT  56.365 155.280 56.645 171.290 ;
        RECT  57.120 155.300 57.400 171.290 ;
        RECT  57.835 155.130 58.115 171.290 ;
        RECT  0.600 155.310 64.400 171.290 ;
        RECT  53.895 155.310 55.870 171.370 ;
        RECT  3.210 155.310 3.490 171.380 ;
        RECT  34.655 155.310 38.715 171.480 ;
        RECT  39.605 155.310 42.020 171.480 ;
        RECT  2.000 0.000 63.000 60.210 ;
        RECT  0.600 0.600 64.400 60.210 ;
        RECT  0.600 0.600 1.210 135.520 ;
        RECT  0.600 91.020 64.400 135.520 ;
        RECT  4.080 91.020 60.940 135.690 ;
        RECT  62.580 91.020 62.995 135.710 ;
        LAYER M3 ;
        RECT  0.600 247.660 23.220 248.740 ;
        RECT  0.600 247.660 22.900 249.400 ;
        RECT  26.260 247.660 64.400 248.740 ;
        RECT  26.580 247.660 27.000 249.400 ;
        RECT  30.440 247.660 64.400 249.400 ;
        RECT  0.600 124.090 64.400 129.850 ;
        RECT  3.990 123.970 60.900 135.790 ;
        RECT  1.640 124.090 63.600 135.790 ;
        RECT  1.810 124.090 2.830 154.520 ;
        RECT  5.155 123.970 60.900 171.560 ;
        RECT  1.640 155.040 63.600 171.560 ;
        RECT  1.640 183.580 63.600 185.950 ;
        RECT  5.490 124.090 63.600 200.820 ;
        RECT  1.640 196.170 63.600 200.820 ;
        RECT  0.600 0.600 64.400 60.480 ;
        RECT  2.000 0.000 63.000 88.700 ;
        RECT  0.600 0.600 1.480 91.220 ;
        RECT  0.600 90.750 64.400 91.220 ;
        LAYER TOP_M ;
        RECT  0.600 247.690 64.400 248.850 ;
        RECT  0.600 247.690 23.010 249.400 ;
        RECT  26.470 247.690 27.110 249.400 ;
        RECT  30.330 247.690 64.400 249.400 ;
        RECT  2.000 0.000 63.000 91.190 ;
        RECT  0.600 0.600 64.400 91.190 ;
    END
END pt3t01d

MACRO pt3t01
    CLASS PAD ;
    FOREIGN pt3t01 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 65.000 BY 250.000 ;
    SYMMETRY X Y R90 ;
    SITE IOSite_c ;
    PIN PAD
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 55.440  LAYER TOP_M  ;
        ANTENNAPARTIALMETALSIDEAREA 287.938  LAYER M3  ;
        ANTENNAPARTIALMETALSIDEAREA 480.740  LAYER M2  ;
        ANTENNADIFFAREA 2657.280  LAYER TOP_M  ;
        ANTENNADIFFAREA 2657.280  LAYER M3  ;
        ANTENNADIFFAREA 1209.600  LAYER M2  ;
        ANTENNAPARTIALCUTAREA 632.318  LAYER TOP_V  ;
        ANTENNAPARTIALCUTAREA 349.898  LAYER V3  ;
        ANTENNAPARTIALCUTAREA 255.798  LAYER V2  ;
        PORT
        LAYER M3 ;
        RECT  23.740 249.580 25.740 250.000 ;
        LAYER M2 ;
        RECT  2.000 61.000 63.000 90.230 ;
        RECT  23.740 246.275 25.740 250.000 ;
        END
    END PAD
    PIN OEN
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 81.726  LAYER M2  ;
        ANTENNAPARTIALMETALSIDEAREA 67.374  LAYER M1  ;
        ANTENNAPARTIALMETALSIDEAREA 41.679  LAYER M3  ;
        ANTENNADIFFAREA 0.250  LAYER M3  ;
        ANTENNAPARTIALCUTAREA 0.203  LAYER V2  ;
        ANTENNAPARTIALCUTAREA 0.135  LAYER V3  ;
        ANTENNAGATEAREA 8.100  LAYER M2  ;
        ANTENNAGATEAREA 9.900  LAYER M3  ;
        PORT
        LAYER M3 ;
        RECT  28.870 249.580 29.600 250.000 ;
        LAYER M2 ;
        RECT  28.870 249.580 29.600 250.000 ;
        END
    END OEN
    PIN I
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 67.374  LAYER M1  ;
        ANTENNAPARTIALMETALSIDEAREA 80.804  LAYER M2  ;
        ANTENNAPARTIALMETALSIDEAREA 41.096  LAYER M3  ;
        ANTENNADIFFAREA 0.250  LAYER M3  ;
        ANTENNAPARTIALCUTAREA 0.203  LAYER V2  ;
        ANTENNAPARTIALCUTAREA 0.135  LAYER V3  ;
        ANTENNAGATEAREA 8.100  LAYER M2  ;
        ANTENNAGATEAREA 9.900  LAYER M3  ;
        PORT
        LAYER M3 ;
        RECT  27.840 249.580 28.570 250.000 ;
        LAYER M2 ;
        RECT  27.840 249.580 28.570 250.000 ;
        END
    END I
    PIN VDDO
        DIRECTION INOUT ;
        USE power ;
        PORT
        LAYER M3 ;
        RECT  64.200 192.330 65.000 200.640 ;
        RECT  0.000 201.660 65.000 221.520 ;
        RECT  0.000 222.720 65.000 246.820 ;
        RECT  0.000 192.330 0.800 200.640 ;
        LAYER M2 ;
        RECT  0.000 186.470 65.000 195.650 ;
        LAYER TOP_M ;
        RECT  0.000 195.170 65.000 200.640 ;
        RECT  0.000 201.660 65.000 221.520 ;
        RECT  0.000 222.720 65.000 246.820 ;
        END
    END VDDO
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        PORT
        LAYER M3 ;
        RECT  64.200 163.510 65.000 190.890 ;
        RECT  0.000 163.510 0.800 190.890 ;
        LAYER M2 ;
        RECT  0.000 172.080 65.000 183.060 ;
        LAYER TOP_M ;
        RECT  0.000 163.500 65.000 194.560 ;
        END
    END VDD
    PIN VSSO
        DIRECTION INOUT ;
        USE ground ;
        PORT
        LAYER M3 ;
        RECT  0.000 92.060 65.000 123.250 ;
        RECT  64.200 149.940 65.000 162.610 ;
        RECT  0.000 149.940 0.800 162.610 ;
        LAYER M2 ;
        RECT  0.000 147.040 65.000 154.520 ;
        LAYER TOP_M ;
        RECT  0.000 92.060 65.000 123.250 ;
        RECT  0.000 155.410 65.000 162.610 ;
        END
    END VSSO
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        PORT
        LAYER M3 ;
        RECT  64.200 130.690 65.000 148.880 ;
        RECT  0.000 130.690 0.800 148.880 ;
        LAYER M2 ;
        RECT  0.000 136.310 65.000 146.340 ;
        LAYER TOP_M ;
        RECT  0.000 123.850 65.000 154.560 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  2.000 0.000 63.000 250.000 ;
        RECT  0.000 88.990 65.000 130.360 ;
        RECT  0.000 136.510 65.000 157.550 ;
        RECT  0.315 158.150 64.700 158.460 ;
        RECT  0.300 158.930 64.700 159.230 ;
        RECT  0.300 159.530 64.700 159.830 ;
        RECT  0.300 160.130 64.700 160.430 ;
        RECT  0.300 160.730 64.700 161.030 ;
        RECT  0.300 161.330 64.700 161.630 ;
        RECT  0.300 161.910 64.700 162.190 ;
        RECT  0.300 162.490 64.700 162.770 ;
        RECT  0.300 163.070 64.700 163.350 ;
        RECT  0.300 163.650 64.700 163.950 ;
        RECT  0.300 164.250 64.700 164.550 ;
        RECT  0.300 164.850 64.700 165.150 ;
        RECT  0.300 165.450 64.700 165.750 ;
        RECT  0.300 166.050 64.700 166.350 ;
        RECT  0.300 166.650 64.700 166.960 ;
        RECT  0.300 167.260 64.700 167.560 ;
        RECT  0.300 167.860 64.700 168.160 ;
        RECT  0.000 169.150 65.000 197.240 ;
        RECT  0.600 0.600 64.400 250.000 ;
        RECT  0.000 198.470 65.000 250.000 ;
        LAYER M2 ;
        RECT  63.180 196.430 63.670 249.400 ;
        RECT  0.600 196.440 64.400 245.485 ;
        RECT  26.530 196.440 64.400 248.790 ;
        RECT  0.600 196.440 22.950 249.400 ;
        RECT  26.530 196.440 27.050 249.400 ;
        RECT  30.390 196.440 64.400 249.400 ;
        RECT  0.600 183.850 64.400 185.680 ;
        RECT  46.230 183.850 51.730 185.870 ;
        RECT  19.790 155.160 20.140 171.290 ;
        RECT  20.440 155.140 20.760 171.290 ;
        RECT  53.655 155.035 53.935 171.290 ;
        RECT  56.365 155.280 56.645 171.290 ;
        RECT  57.120 155.300 57.400 171.290 ;
        RECT  57.835 155.130 58.115 171.290 ;
        RECT  0.600 155.310 64.400 171.290 ;
        RECT  53.895 155.310 55.870 171.370 ;
        RECT  3.210 155.310 3.490 171.380 ;
        RECT  34.655 155.310 38.715 171.480 ;
        RECT  39.605 155.310 42.020 171.480 ;
        RECT  2.000 0.000 63.000 60.210 ;
        RECT  0.600 0.600 64.400 60.210 ;
        RECT  0.600 0.600 1.210 135.520 ;
        RECT  0.600 91.020 64.400 135.520 ;
        RECT  4.080 91.020 60.940 135.690 ;
        RECT  62.580 91.020 62.995 135.710 ;
        LAYER M3 ;
        RECT  0.600 247.660 23.220 248.740 ;
        RECT  0.600 247.660 22.900 249.400 ;
        RECT  26.260 247.660 64.400 248.740 ;
        RECT  26.580 247.660 27.000 249.400 ;
        RECT  30.440 247.660 64.400 249.400 ;
        RECT  0.600 124.090 64.400 129.850 ;
        RECT  3.990 123.970 60.900 135.790 ;
        RECT  1.640 124.090 63.600 135.790 ;
        RECT  1.810 124.090 2.830 154.520 ;
        RECT  5.155 123.970 60.900 171.560 ;
        RECT  1.640 155.040 63.600 171.560 ;
        RECT  1.640 183.580 63.600 185.950 ;
        RECT  5.490 124.090 63.600 200.820 ;
        RECT  1.640 196.170 63.600 200.820 ;
        RECT  0.600 0.600 64.400 60.480 ;
        RECT  2.000 0.000 63.000 88.700 ;
        RECT  0.600 0.600 1.480 91.220 ;
        RECT  0.600 90.750 64.400 91.220 ;
        LAYER TOP_M ;
        RECT  0.600 247.690 64.400 248.850 ;
        RECT  0.600 247.690 23.010 249.400 ;
        RECT  26.470 247.690 27.110 249.400 ;
        RECT  30.330 247.690 64.400 249.400 ;
        RECT  2.000 0.000 63.000 91.190 ;
        RECT  0.600 0.600 64.400 91.190 ;
    END
END pt3t01

MACRO pt3o03
    CLASS PAD ;
    FOREIGN pt3o03 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 65.000 BY 250.000 ;
    SYMMETRY X Y R90 ;
    SITE IOSite_c ;
    PIN PAD
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 55.440  LAYER TOP_M  ;
        ANTENNAPARTIALMETALSIDEAREA 287.938  LAYER M3  ;
        ANTENNAPARTIALMETALSIDEAREA 480.740  LAYER M2  ;
        ANTENNADIFFAREA 2657.280  LAYER TOP_M  ;
        ANTENNADIFFAREA 2657.280  LAYER M3  ;
        ANTENNADIFFAREA 1209.600  LAYER M2  ;
        ANTENNAPARTIALCUTAREA 632.318  LAYER TOP_V  ;
        ANTENNAPARTIALCUTAREA 349.898  LAYER V3  ;
        ANTENNAPARTIALCUTAREA 255.798  LAYER V2  ;
        PORT
        LAYER M3 ;
        RECT  26.310 249.580 28.310 250.000 ;
        LAYER M2 ;
        RECT  2.000 61.000 63.000 90.230 ;
        RECT  26.310 246.275 28.310 250.000 ;
        END
    END PAD
    PIN I
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 67.374  LAYER M1  ;
        ANTENNAPARTIALMETALSIDEAREA 81.652  LAYER M2  ;
        ANTENNAPARTIALMETALSIDEAREA 41.425  LAYER M3  ;
        ANTENNADIFFAREA 0.250  LAYER M3  ;
        ANTENNAPARTIALCUTAREA 0.338  LAYER V2  ;
        ANTENNAPARTIALCUTAREA 0.135  LAYER V3  ;
        ANTENNAGATEAREA 18.900  LAYER M2  ;
        ANTENNAGATEAREA 20.700  LAYER M3  ;
        PORT
        LAYER M3 ;
        RECT  30.310 249.580 31.040 250.000 ;
        LAYER M2 ;
        RECT  30.310 249.580 31.040 250.000 ;
        END
    END I
    PIN VDDO
        DIRECTION INOUT ;
        USE power ;
        PORT
        LAYER M3 ;
        RECT  64.200 192.330 65.000 200.640 ;
        RECT  0.000 201.660 65.000 221.520 ;
        RECT  0.000 222.720 65.000 246.820 ;
        RECT  0.000 192.330 0.800 200.640 ;
        LAYER M2 ;
        RECT  0.000 186.470 65.000 195.650 ;
        LAYER TOP_M ;
        RECT  0.000 195.170 65.000 200.640 ;
        RECT  0.000 201.660 65.000 221.520 ;
        RECT  0.000 222.720 65.000 246.820 ;
        END
    END VDDO
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        PORT
        LAYER M3 ;
        RECT  64.200 163.510 65.000 190.890 ;
        RECT  0.000 163.510 0.800 190.890 ;
        LAYER M2 ;
        RECT  0.000 172.080 65.000 183.060 ;
        LAYER TOP_M ;
        RECT  0.000 163.500 65.000 194.560 ;
        END
    END VDD
    PIN VSSO
        DIRECTION INOUT ;
        USE ground ;
        PORT
        LAYER M3 ;
        RECT  0.000 92.060 65.000 123.250 ;
        RECT  64.200 149.940 65.000 162.610 ;
        RECT  0.000 149.940 0.800 162.610 ;
        LAYER M2 ;
        RECT  0.000 147.040 65.000 154.520 ;
        LAYER TOP_M ;
        RECT  0.000 92.060 65.000 123.250 ;
        RECT  0.000 155.410 65.000 162.610 ;
        END
    END VSSO
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        PORT
        LAYER M3 ;
        RECT  64.200 130.690 65.000 148.880 ;
        RECT  0.000 130.690 0.800 148.880 ;
        LAYER M2 ;
        RECT  0.000 136.310 65.000 146.340 ;
        LAYER TOP_M ;
        RECT  0.000 123.850 65.000 154.560 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  2.000 0.000 63.000 250.000 ;
        RECT  0.000 88.990 65.000 130.360 ;
        RECT  0.000 136.510 65.000 157.550 ;
        RECT  0.300 158.930 64.700 159.230 ;
        RECT  0.300 159.530 64.700 159.830 ;
        RECT  0.300 160.130 64.700 160.430 ;
        RECT  0.300 160.730 64.700 161.030 ;
        RECT  0.300 161.330 64.700 161.630 ;
        RECT  0.300 161.910 64.700 162.190 ;
        RECT  0.300 162.490 64.700 162.770 ;
        RECT  0.300 163.070 64.700 163.350 ;
        RECT  0.300 163.650 64.700 163.950 ;
        RECT  0.300 164.250 64.700 164.550 ;
        RECT  0.300 164.850 64.700 165.150 ;
        RECT  0.300 165.450 64.700 165.750 ;
        RECT  0.300 166.050 64.700 166.350 ;
        RECT  0.300 166.650 64.700 166.960 ;
        RECT  0.300 167.260 64.700 167.560 ;
        RECT  0.300 167.860 64.700 168.160 ;
        RECT  0.000 169.150 65.000 197.240 ;
        RECT  0.600 0.600 64.400 250.000 ;
        RECT  0.000 198.470 65.000 250.000 ;
        LAYER M2 ;
        RECT  2.800 196.110 3.220 249.400 ;
        RECT  63.180 196.430 63.670 249.400 ;
        RECT  0.600 196.440 64.400 245.485 ;
        RECT  29.100 196.440 64.400 248.790 ;
        RECT  0.600 196.440 25.520 249.400 ;
        RECT  29.100 196.440 29.520 249.400 ;
        RECT  31.830 196.440 64.400 249.400 ;
        RECT  55.890 183.790 56.190 185.680 ;
        RECT  58.060 183.750 58.350 185.680 ;
        RECT  0.600 183.850 64.400 185.680 ;
        RECT  46.070 183.850 51.600 185.820 ;
        RECT  8.170 155.125 8.490 171.290 ;
        RECT  43.245 155.035 43.525 171.290 ;
        RECT  45.955 155.280 46.235 171.370 ;
        RECT  47.425 155.130 47.705 171.370 ;
        RECT  58.295 155.175 58.605 171.290 ;
        RECT  60.755 155.175 61.065 171.290 ;
        RECT  63.290 155.270 63.600 171.290 ;
        RECT  0.600 155.310 64.400 171.290 ;
        RECT  43.485 155.310 56.355 171.370 ;
        RECT  29.195 155.310 31.610 171.480 ;
        RECT  2.000 0.000 63.000 60.210 ;
        RECT  0.600 0.600 64.400 60.210 ;
        RECT  0.600 0.600 1.210 135.520 ;
        RECT  0.600 91.020 64.400 135.520 ;
        RECT  4.080 91.020 60.940 135.690 ;
        LAYER M3 ;
        RECT  0.600 247.660 25.790 248.740 ;
        RECT  0.600 247.660 25.470 249.400 ;
        RECT  28.830 247.660 64.400 248.740 ;
        RECT  29.150 247.660 29.470 249.400 ;
        RECT  31.880 247.660 64.400 249.400 ;
        RECT  4.040 123.850 60.900 200.820 ;
        RECT  0.600 124.090 64.400 129.850 ;
        RECT  1.640 124.090 63.600 135.790 ;
        RECT  1.810 124.090 2.830 154.520 ;
        RECT  1.640 155.040 63.600 171.560 ;
        RECT  1.640 183.580 63.600 185.950 ;
        RECT  2.800 155.040 63.600 200.820 ;
        RECT  3.340 124.090 63.600 200.820 ;
        RECT  1.640 196.170 63.600 200.820 ;
        RECT  0.600 0.600 64.400 60.480 ;
        RECT  2.000 0.000 63.000 88.700 ;
        RECT  0.600 0.600 1.480 91.220 ;
        RECT  0.600 90.750 64.400 91.220 ;
        LAYER TOP_M ;
        RECT  0.600 247.690 64.400 248.850 ;
        RECT  0.600 247.690 25.580 249.400 ;
        RECT  29.040 247.690 29.580 249.400 ;
        RECT  31.770 247.690 64.400 249.400 ;
        RECT  2.000 0.000 63.000 91.190 ;
        RECT  0.600 0.600 64.400 91.190 ;
    END
END pt3o03

MACRO pt3o02
    CLASS PAD ;
    FOREIGN pt3o02 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 65.000 BY 250.000 ;
    SYMMETRY X Y R90 ;
    SITE IOSite_c ;
    PIN PAD
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 55.440  LAYER TOP_M  ;
        ANTENNAPARTIALMETALSIDEAREA 287.938  LAYER M3  ;
        ANTENNAPARTIALMETALSIDEAREA 480.740  LAYER M2  ;
        ANTENNADIFFAREA 2657.280  LAYER TOP_M  ;
        ANTENNADIFFAREA 2657.280  LAYER M3  ;
        ANTENNADIFFAREA 1209.600  LAYER M2  ;
        ANTENNAPARTIALCUTAREA 632.318  LAYER TOP_V  ;
        ANTENNAPARTIALCUTAREA 349.898  LAYER V3  ;
        ANTENNAPARTIALCUTAREA 255.798  LAYER V2  ;
        PORT
        LAYER M3 ;
        RECT  26.310 249.580 28.310 250.000 ;
        LAYER M2 ;
        RECT  2.000 61.000 63.000 90.230 ;
        RECT  26.310 246.275 28.310 250.000 ;
        END
    END PAD
    PIN I
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 67.374  LAYER M1  ;
        ANTENNAPARTIALMETALSIDEAREA 81.652  LAYER M2  ;
        ANTENNAPARTIALMETALSIDEAREA 41.425  LAYER M3  ;
        ANTENNADIFFAREA 0.250  LAYER M3  ;
        ANTENNAPARTIALCUTAREA 0.338  LAYER V2  ;
        ANTENNAPARTIALCUTAREA 0.135  LAYER V3  ;
        ANTENNAGATEAREA 18.900  LAYER M2  ;
        ANTENNAGATEAREA 20.700  LAYER M3  ;
        PORT
        LAYER M3 ;
        RECT  30.310 249.580 31.040 250.000 ;
        LAYER M2 ;
        RECT  30.310 249.580 31.040 250.000 ;
        END
    END I
    PIN VDDO
        DIRECTION INOUT ;
        USE power ;
        PORT
        LAYER M3 ;
        RECT  64.200 192.330 65.000 200.640 ;
        RECT  0.000 201.660 65.000 221.520 ;
        RECT  0.000 222.720 65.000 246.820 ;
        RECT  0.000 192.330 0.800 200.640 ;
        LAYER M2 ;
        RECT  0.000 186.470 65.000 195.650 ;
        LAYER TOP_M ;
        RECT  0.000 195.170 65.000 200.640 ;
        RECT  0.000 201.660 65.000 221.520 ;
        RECT  0.000 222.720 65.000 246.820 ;
        END
    END VDDO
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        PORT
        LAYER M3 ;
        RECT  64.200 163.510 65.000 190.890 ;
        RECT  0.000 163.510 0.800 190.890 ;
        LAYER M2 ;
        RECT  0.000 172.080 65.000 183.060 ;
        LAYER TOP_M ;
        RECT  0.000 163.500 65.000 194.560 ;
        END
    END VDD
    PIN VSSO
        DIRECTION INOUT ;
        USE ground ;
        PORT
        LAYER M3 ;
        RECT  0.000 92.060 65.000 123.250 ;
        RECT  64.200 149.940 65.000 162.610 ;
        RECT  0.000 149.940 0.800 162.610 ;
        LAYER M2 ;
        RECT  0.000 147.040 65.000 154.520 ;
        LAYER TOP_M ;
        RECT  0.000 92.060 65.000 123.250 ;
        RECT  0.000 155.410 65.000 162.610 ;
        END
    END VSSO
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        PORT
        LAYER M3 ;
        RECT  64.200 130.690 65.000 148.880 ;
        RECT  0.000 130.690 0.800 148.880 ;
        LAYER M2 ;
        RECT  0.000 136.310 65.000 146.340 ;
        LAYER TOP_M ;
        RECT  0.000 123.850 65.000 154.560 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  2.000 0.000 63.000 250.000 ;
        RECT  0.000 88.990 65.000 130.360 ;
        RECT  0.000 136.510 65.000 157.550 ;
        RECT  0.300 158.930 64.700 159.230 ;
        RECT  0.300 159.530 64.700 159.830 ;
        RECT  0.300 160.130 64.700 160.430 ;
        RECT  0.300 160.730 64.700 161.030 ;
        RECT  0.300 161.330 64.700 161.630 ;
        RECT  0.300 161.910 64.700 162.190 ;
        RECT  0.300 162.490 64.700 162.770 ;
        RECT  0.300 163.070 64.700 163.350 ;
        RECT  0.300 163.650 64.700 163.950 ;
        RECT  0.300 164.250 64.700 164.550 ;
        RECT  0.300 164.850 64.700 165.150 ;
        RECT  0.300 165.450 64.700 165.750 ;
        RECT  0.300 166.050 64.700 166.350 ;
        RECT  0.300 166.650 64.700 166.960 ;
        RECT  0.300 167.260 64.700 167.560 ;
        RECT  0.300 167.860 64.700 168.160 ;
        RECT  0.000 169.150 65.000 197.240 ;
        RECT  0.600 0.600 64.400 250.000 ;
        RECT  0.000 198.470 65.000 250.000 ;
        LAYER M2 ;
        RECT  2.800 196.110 3.220 249.400 ;
        RECT  63.180 196.430 63.670 249.400 ;
        RECT  0.600 196.440 64.400 245.485 ;
        RECT  29.100 196.440 64.400 248.790 ;
        RECT  0.600 196.440 25.520 249.400 ;
        RECT  29.100 196.440 29.520 249.400 ;
        RECT  31.830 196.440 64.400 249.400 ;
        RECT  55.890 183.790 56.190 185.680 ;
        RECT  58.060 183.750 58.350 185.680 ;
        RECT  0.600 183.850 64.400 185.680 ;
        RECT  46.070 183.850 51.600 185.820 ;
        RECT  8.170 155.125 8.490 171.290 ;
        RECT  43.245 155.035 43.525 171.290 ;
        RECT  45.955 155.280 46.235 171.370 ;
        RECT  47.425 155.130 47.705 171.370 ;
        RECT  58.045 155.175 58.355 171.290 ;
        RECT  60.505 155.175 60.815 171.290 ;
        RECT  63.040 155.270 63.350 171.290 ;
        RECT  0.600 155.310 64.400 171.290 ;
        RECT  43.485 155.310 56.355 171.370 ;
        RECT  29.195 155.310 31.610 171.480 ;
        RECT  2.000 0.000 63.000 60.210 ;
        RECT  0.600 0.600 64.400 60.210 ;
        RECT  0.600 0.600 1.210 135.520 ;
        RECT  0.600 91.020 64.400 135.520 ;
        RECT  4.080 91.020 60.940 135.690 ;
        LAYER M3 ;
        RECT  0.600 247.660 25.790 248.740 ;
        RECT  0.600 247.660 25.470 249.400 ;
        RECT  28.830 247.660 64.400 248.740 ;
        RECT  29.150 247.660 29.470 249.400 ;
        RECT  31.880 247.660 64.400 249.400 ;
        RECT  4.040 123.970 60.900 200.820 ;
        RECT  0.600 124.090 64.400 129.850 ;
        RECT  1.640 124.090 63.600 135.790 ;
        RECT  1.810 124.090 2.830 154.520 ;
        RECT  1.640 155.040 63.600 171.560 ;
        RECT  1.640 183.580 63.600 185.950 ;
        RECT  2.800 155.040 63.600 200.820 ;
        RECT  3.230 124.090 63.600 200.820 ;
        RECT  1.640 196.170 63.600 200.820 ;
        RECT  0.600 0.600 64.400 60.480 ;
        RECT  2.000 0.000 63.000 88.700 ;
        RECT  0.600 0.600 1.480 91.220 ;
        RECT  0.600 90.750 64.400 91.220 ;
        LAYER TOP_M ;
        RECT  0.600 247.690 64.400 248.850 ;
        RECT  0.600 247.690 25.580 249.400 ;
        RECT  29.040 247.690 29.580 249.400 ;
        RECT  31.770 247.690 64.400 249.400 ;
        RECT  2.000 0.000 63.000 91.190 ;
        RECT  0.600 0.600 64.400 91.190 ;
    END
END pt3o02

MACRO pt3o01
    CLASS PAD ;
    FOREIGN pt3o01 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 65.000 BY 250.000 ;
    SYMMETRY X Y R90 ;
    SITE IOSite_c ;
    PIN PAD
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 55.440  LAYER TOP_M  ;
        ANTENNAPARTIALMETALSIDEAREA 287.938  LAYER M3  ;
        ANTENNAPARTIALMETALSIDEAREA 480.740  LAYER M2  ;
        ANTENNADIFFAREA 2657.280  LAYER TOP_M  ;
        ANTENNADIFFAREA 2657.280  LAYER M3  ;
        ANTENNADIFFAREA 1209.600  LAYER M2  ;
        ANTENNAPARTIALCUTAREA 632.318  LAYER TOP_V  ;
        ANTENNAPARTIALCUTAREA 349.898  LAYER V3  ;
        ANTENNAPARTIALCUTAREA 255.798  LAYER V2  ;
        PORT
        LAYER M3 ;
        RECT  26.310 249.580 28.310 250.000 ;
        LAYER M2 ;
        RECT  2.000 61.000 63.000 90.230 ;
        RECT  26.310 246.275 28.310 250.000 ;
        END
    END PAD
    PIN I
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 67.374  LAYER M1  ;
        ANTENNAPARTIALMETALSIDEAREA 81.652  LAYER M2  ;
        ANTENNAPARTIALMETALSIDEAREA 41.425  LAYER M3  ;
        ANTENNADIFFAREA 0.250  LAYER M3  ;
        ANTENNAPARTIALCUTAREA 0.135  LAYER V3  ;
        ANTENNAPARTIALCUTAREA 0.270  LAYER V2  ;
        ANTENNAGATEAREA 8.100  LAYER M2  ;
        ANTENNAGATEAREA 9.900  LAYER M3  ;
        PORT
        LAYER M3 ;
        RECT  30.310 249.580 31.040 250.000 ;
        LAYER M2 ;
        RECT  30.310 249.580 31.040 250.000 ;
        END
    END I
    PIN VDDO
        DIRECTION INOUT ;
        USE power ;
        PORT
        LAYER M3 ;
        RECT  64.200 192.330 65.000 200.640 ;
        RECT  0.000 201.660 65.000 221.520 ;
        RECT  0.000 222.720 65.000 246.820 ;
        RECT  0.000 192.330 0.800 200.640 ;
        LAYER M2 ;
        RECT  0.000 186.470 65.000 195.650 ;
        LAYER TOP_M ;
        RECT  0.000 195.170 65.000 200.640 ;
        RECT  0.000 201.660 65.000 221.520 ;
        RECT  0.000 222.720 65.000 246.820 ;
        END
    END VDDO
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        PORT
        LAYER M3 ;
        RECT  64.200 163.510 65.000 190.890 ;
        RECT  0.000 163.510 0.800 190.890 ;
        LAYER M2 ;
        RECT  0.000 172.080 65.000 183.060 ;
        LAYER TOP_M ;
        RECT  0.000 163.500 65.000 194.560 ;
        END
    END VDD
    PIN VSSO
        DIRECTION INOUT ;
        USE ground ;
        PORT
        LAYER M3 ;
        RECT  0.000 92.060 65.000 123.250 ;
        RECT  64.200 149.940 65.000 162.610 ;
        RECT  0.000 149.940 0.800 162.610 ;
        LAYER M2 ;
        RECT  0.000 147.040 65.000 154.520 ;
        LAYER TOP_M ;
        RECT  0.000 92.060 65.000 123.250 ;
        RECT  0.000 155.410 65.000 162.610 ;
        END
    END VSSO
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        PORT
        LAYER M3 ;
        RECT  64.200 130.690 65.000 148.880 ;
        RECT  0.000 130.690 0.800 148.880 ;
        LAYER M2 ;
        RECT  0.000 136.310 65.000 146.340 ;
        LAYER TOP_M ;
        RECT  0.000 123.850 65.000 154.560 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  2.000 0.000 63.000 250.000 ;
        RECT  0.000 88.990 65.000 130.360 ;
        RECT  0.000 136.510 65.000 157.550 ;
        RECT  0.300 158.930 64.700 159.230 ;
        RECT  0.300 159.530 64.700 159.830 ;
        RECT  0.300 160.130 64.700 160.430 ;
        RECT  0.300 160.730 64.700 161.030 ;
        RECT  0.300 161.330 64.700 161.630 ;
        RECT  0.300 161.910 64.700 162.190 ;
        RECT  0.300 162.490 64.700 162.770 ;
        RECT  0.300 163.070 64.700 163.350 ;
        RECT  0.300 163.650 64.700 163.950 ;
        RECT  0.300 164.250 64.700 164.550 ;
        RECT  0.300 164.850 64.700 165.150 ;
        RECT  0.300 165.450 64.700 165.750 ;
        RECT  0.300 166.050 64.700 166.350 ;
        RECT  0.300 166.650 64.700 166.960 ;
        RECT  0.300 167.260 64.700 167.560 ;
        RECT  0.300 167.860 64.700 168.160 ;
        RECT  0.000 169.150 65.000 197.240 ;
        RECT  0.600 0.600 64.400 250.000 ;
        RECT  0.000 198.470 65.000 250.000 ;
        LAYER M2 ;
        RECT  2.520 196.270 2.940 249.400 ;
        RECT  63.180 196.430 63.670 249.400 ;
        RECT  0.600 196.440 64.400 245.485 ;
        RECT  29.100 196.440 64.400 248.790 ;
        RECT  0.600 196.440 25.520 249.400 ;
        RECT  29.100 196.440 29.520 249.400 ;
        RECT  31.830 196.440 64.400 249.400 ;
        RECT  55.890 183.790 56.190 185.680 ;
        RECT  58.060 183.750 58.350 185.680 ;
        RECT  0.600 183.850 64.400 185.680 ;
        RECT  46.070 183.850 51.600 185.820 ;
        RECT  43.245 155.035 43.525 171.290 ;
        RECT  45.955 155.280 46.235 171.370 ;
        RECT  47.425 155.130 47.705 171.370 ;
        RECT  60.705 155.175 61.015 171.290 ;
        RECT  63.290 155.270 63.600 171.290 ;
        RECT  0.600 155.310 64.400 171.290 ;
        RECT  43.485 155.310 56.355 171.370 ;
        RECT  29.195 155.310 31.610 171.480 ;
        RECT  2.000 0.000 63.000 60.210 ;
        RECT  0.600 0.600 64.400 60.210 ;
        RECT  0.600 0.600 1.210 135.520 ;
        RECT  0.600 91.020 64.400 135.520 ;
        RECT  4.080 91.020 60.940 135.690 ;
        LAYER M3 ;
        RECT  0.600 247.660 25.790 248.740 ;
        RECT  0.600 247.660 25.470 249.400 ;
        RECT  28.830 247.660 64.400 248.740 ;
        RECT  29.150 247.660 29.470 249.400 ;
        RECT  31.880 247.660 64.400 249.400 ;
        RECT  4.040 123.870 60.900 200.820 ;
        RECT  0.600 124.090 64.400 129.850 ;
        RECT  1.640 124.090 63.600 135.790 ;
        RECT  1.810 124.090 2.830 154.520 ;
        RECT  1.640 155.040 63.600 171.560 ;
        RECT  1.640 183.580 63.600 185.950 ;
        RECT  2.520 155.040 63.600 200.820 ;
        RECT  4.040 124.090 63.600 200.820 ;
        RECT  1.640 196.170 63.600 200.820 ;
        RECT  0.600 0.600 64.400 60.480 ;
        RECT  2.000 0.000 63.000 88.700 ;
        RECT  0.600 0.600 1.480 91.220 ;
        RECT  0.600 90.750 64.400 91.220 ;
        LAYER TOP_M ;
        RECT  0.600 247.690 64.400 248.850 ;
        RECT  0.600 247.690 25.580 249.400 ;
        RECT  29.040 247.690 29.580 249.400 ;
        RECT  31.770 247.690 64.400 249.400 ;
        RECT  2.000 0.000 63.000 91.190 ;
        RECT  0.600 0.600 64.400 91.190 ;
    END
END pt3o01

MACRO pt3b03u
    CLASS PAD ;
    FOREIGN pt3b03u 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 65.000 BY 250.000 ;
    SYMMETRY X Y R90 ;
    SITE IOSite_c ;
    PIN PAD
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 55.440  LAYER TOP_M  ;
        ANTENNAPARTIALMETALSIDEAREA 287.938  LAYER M3  ;
        ANTENNAPARTIALMETALSIDEAREA 480.740  LAYER M2  ;
        ANTENNADIFFAREA 2657.280  LAYER TOP_M  ;
        ANTENNADIFFAREA 2657.280  LAYER M3  ;
        ANTENNADIFFAREA 1209.600  LAYER M2  ;
        ANTENNAPARTIALCUTAREA 632.318  LAYER TOP_V  ;
        ANTENNAPARTIALCUTAREA 349.898  LAYER V3  ;
        ANTENNAPARTIALCUTAREA 255.798  LAYER V2  ;
        PORT
        LAYER M3 ;
        RECT  23.740 249.580 25.740 250.000 ;
        LAYER M2 ;
        RECT  2.000 61.000 63.000 90.230 ;
        RECT  23.740 246.275 25.740 250.000 ;
        END
    END PAD
    PIN CIN
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 32.277  LAYER M3  ;
        ANTENNAPARTIALMETALSIDEAREA 96.916  LAYER M2  ;
        ANTENNAPARTIALMETALSIDEAREA 67.374  LAYER M1  ;
        ANTENNADIFFAREA 20.600  LAYER M3  ;
        ANTENNAPARTIALCUTAREA 0.135  LAYER V3  ;
        ANTENNAPARTIALCUTAREA 0.203  LAYER V2  ;
        PORT
        LAYER M3 ;
        RECT  28.870 249.580 29.600 250.000 ;
        LAYER M2 ;
        RECT  28.870 249.580 29.600 250.000 ;
        END
    END CIN
    PIN OEN
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 80.634  LAYER M2  ;
        ANTENNAPARTIALMETALSIDEAREA 67.374  LAYER M1  ;
        ANTENNAPARTIALMETALSIDEAREA 41.679  LAYER M3  ;
        ANTENNADIFFAREA 0.250  LAYER M3  ;
        ANTENNAPARTIALCUTAREA 0.203  LAYER V2  ;
        ANTENNAPARTIALCUTAREA 0.135  LAYER V3  ;
        ANTENNAGATEAREA 8.100  LAYER M2  ;
        ANTENNAGATEAREA 9.900  LAYER M3  ;
        PORT
        LAYER M3 ;
        RECT  29.900 249.580 30.630 250.000 ;
        LAYER M2 ;
        RECT  29.900 249.580 30.630 250.000 ;
        END
    END OEN
    PIN I
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 67.374  LAYER M1  ;
        ANTENNAPARTIALMETALSIDEAREA 80.804  LAYER M2  ;
        ANTENNAPARTIALMETALSIDEAREA 41.096  LAYER M3  ;
        ANTENNADIFFAREA 0.250  LAYER M3  ;
        ANTENNAPARTIALCUTAREA 0.270  LAYER V2  ;
        ANTENNAPARTIALCUTAREA 0.135  LAYER V3  ;
        ANTENNAGATEAREA 18.900  LAYER M2  ;
        ANTENNAGATEAREA 20.700  LAYER M3  ;
        PORT
        LAYER M3 ;
        RECT  27.840 249.580 28.570 250.000 ;
        LAYER M2 ;
        RECT  27.840 249.580 28.570 250.000 ;
        END
    END I
    PIN VDDO
        DIRECTION INOUT ;
        USE power ;
        PORT
        LAYER M3 ;
        RECT  64.200 192.330 65.000 200.640 ;
        RECT  0.000 201.660 65.000 221.520 ;
        RECT  0.000 222.720 65.000 246.820 ;
        RECT  0.000 192.330 0.800 200.640 ;
        LAYER M2 ;
        RECT  0.000 186.470 65.000 195.650 ;
        LAYER TOP_M ;
        RECT  0.000 195.170 65.000 200.640 ;
        RECT  0.000 201.660 65.000 221.520 ;
        RECT  0.000 222.720 65.000 246.820 ;
        END
    END VDDO
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        PORT
        LAYER M3 ;
        RECT  64.200 163.510 65.000 190.890 ;
        RECT  0.000 163.510 0.800 190.890 ;
        LAYER M2 ;
        RECT  0.000 172.080 65.000 183.060 ;
        LAYER TOP_M ;
        RECT  0.000 163.500 65.000 194.560 ;
        END
    END VDD
    PIN VSSO
        DIRECTION INOUT ;
        USE ground ;
        PORT
        LAYER M3 ;
        RECT  0.000 92.060 65.000 123.250 ;
        RECT  64.200 149.940 65.000 162.610 ;
        RECT  0.000 149.940 0.800 162.610 ;
        LAYER M2 ;
        RECT  0.000 147.040 65.000 154.520 ;
        LAYER TOP_M ;
        RECT  0.000 92.060 65.000 123.250 ;
        RECT  0.000 155.410 65.000 162.610 ;
        END
    END VSSO
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        PORT
        LAYER M3 ;
        RECT  64.200 130.690 65.000 148.880 ;
        RECT  0.000 130.690 0.800 148.880 ;
        LAYER M2 ;
        RECT  0.000 136.310 65.000 146.340 ;
        LAYER TOP_M ;
        RECT  0.000 123.850 65.000 154.560 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  2.000 0.000 63.000 250.000 ;
        RECT  0.000 88.990 65.000 130.360 ;
        RECT  0.000 136.510 65.000 157.550 ;
        RECT  0.315 158.150 64.700 158.460 ;
        RECT  0.300 158.930 64.700 159.230 ;
        RECT  0.300 159.530 64.700 159.830 ;
        RECT  0.300 160.130 64.700 160.430 ;
        RECT  0.300 160.730 64.700 161.030 ;
        RECT  0.300 161.330 64.700 161.630 ;
        RECT  0.300 161.910 64.700 162.190 ;
        RECT  0.300 162.490 64.700 162.770 ;
        RECT  0.300 163.070 64.700 163.350 ;
        RECT  0.300 163.650 64.700 163.950 ;
        RECT  0.300 164.250 64.700 164.550 ;
        RECT  0.300 164.850 64.700 165.150 ;
        RECT  0.300 165.450 64.700 165.750 ;
        RECT  0.300 166.050 64.700 166.350 ;
        RECT  0.300 166.650 64.700 166.960 ;
        RECT  0.300 167.260 64.700 167.560 ;
        RECT  0.300 167.860 64.700 168.160 ;
        RECT  0.000 169.150 65.000 197.240 ;
        RECT  0.600 0.600 64.400 250.000 ;
        RECT  0.000 198.470 65.000 250.000 ;
        LAYER M2 ;
        RECT  1.840 196.420 2.120 249.400 ;
        RECT  63.180 196.430 63.670 249.400 ;
        RECT  0.600 196.440 64.400 245.485 ;
        RECT  26.530 196.440 64.400 248.790 ;
        RECT  0.600 196.440 22.950 249.400 ;
        RECT  26.530 196.440 27.050 249.400 ;
        RECT  31.420 196.440 64.400 249.400 ;
        RECT  19.440 183.720 52.225 185.680 ;
        RECT  0.600 183.850 64.400 185.680 ;
        RECT  46.230 183.720 51.730 185.870 ;
        RECT  55.235 183.850 56.645 185.900 ;
        RECT  4.480 154.920 7.530 171.290 ;
        RECT  8.170 155.125 8.490 171.290 ;
        RECT  22.160 155.160 22.510 171.290 ;
        RECT  22.810 155.140 23.130 171.290 ;
        RECT  31.960 155.120 35.830 171.290 ;
        RECT  53.655 155.035 53.935 171.290 ;
        RECT  56.365 155.280 56.645 171.315 ;
        RECT  57.120 155.300 57.400 171.315 ;
        RECT  57.835 155.130 58.115 171.315 ;
        RECT  0.600 155.310 64.400 171.290 ;
        RECT  56.240 155.310 61.880 171.315 ;
        RECT  53.895 155.310 55.870 171.370 ;
        RECT  3.170 155.310 3.450 171.380 ;
        RECT  34.655 155.310 38.715 171.480 ;
        RECT  39.605 155.310 42.020 171.480 ;
        RECT  2.000 0.000 63.000 60.210 ;
        RECT  0.600 0.600 64.400 60.210 ;
        RECT  0.600 0.600 1.210 135.520 ;
        RECT  0.600 91.020 64.400 135.520 ;
        RECT  4.080 91.020 60.940 135.690 ;
        RECT  62.580 91.020 62.995 135.710 ;
        LAYER M3 ;
        RECT  0.600 247.660 23.220 248.740 ;
        RECT  0.600 247.660 22.900 249.400 ;
        RECT  26.260 247.660 64.400 248.740 ;
        RECT  26.580 247.660 27.000 249.400 ;
        RECT  31.470 247.660 64.400 249.400 ;
        RECT  0.600 124.090 64.400 129.850 ;
        RECT  1.640 124.090 63.600 135.790 ;
        RECT  1.810 124.090 2.830 154.520 ;
        RECT  3.510 124.090 63.600 171.560 ;
        RECT  4.040 123.970 60.900 171.560 ;
        RECT  1.640 155.040 63.600 171.560 ;
        RECT  1.640 183.580 63.600 185.950 ;
        RECT  5.515 124.090 63.600 200.820 ;
        RECT  1.640 196.170 63.600 200.820 ;
        RECT  56.300 123.970 56.580 201.060 ;
        RECT  0.600 0.600 64.400 60.480 ;
        RECT  2.000 0.000 63.000 88.700 ;
        RECT  0.600 0.600 1.480 91.220 ;
        RECT  0.600 90.750 64.400 91.220 ;
        LAYER TOP_M ;
        RECT  0.600 247.690 64.400 248.850 ;
        RECT  0.600 247.690 23.010 249.400 ;
        RECT  26.470 247.690 27.110 249.400 ;
        RECT  31.360 247.690 64.400 249.400 ;
        RECT  2.000 0.000 63.000 91.190 ;
        RECT  0.600 0.600 64.400 91.190 ;
    END
END pt3b03u

MACRO pt3b03d
    CLASS PAD ;
    FOREIGN pt3b03d 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 65.000 BY 250.000 ;
    SYMMETRY X Y R90 ;
    SITE IOSite_c ;
    PIN PAD
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 55.440  LAYER TOP_M  ;
        ANTENNAPARTIALMETALSIDEAREA 287.938  LAYER M3  ;
        ANTENNAPARTIALMETALSIDEAREA 480.740  LAYER M2  ;
        ANTENNADIFFAREA 2657.280  LAYER TOP_M  ;
        ANTENNADIFFAREA 2657.280  LAYER M3  ;
        ANTENNADIFFAREA 1209.600  LAYER M2  ;
        ANTENNAPARTIALCUTAREA 632.318  LAYER TOP_V  ;
        ANTENNAPARTIALCUTAREA 349.898  LAYER V3  ;
        ANTENNAPARTIALCUTAREA 255.798  LAYER V2  ;
        PORT
        LAYER M3 ;
        RECT  23.740 249.580 25.740 250.000 ;
        LAYER M2 ;
        RECT  2.000 61.000 63.000 90.230 ;
        RECT  23.740 246.275 25.740 250.000 ;
        END
    END PAD
    PIN CIN
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 32.277  LAYER M3  ;
        ANTENNAPARTIALMETALSIDEAREA 96.916  LAYER M2  ;
        ANTENNAPARTIALMETALSIDEAREA 67.374  LAYER M1  ;
        ANTENNADIFFAREA 20.600  LAYER M3  ;
        ANTENNAPARTIALCUTAREA 0.135  LAYER V3  ;
        ANTENNAPARTIALCUTAREA 0.203  LAYER V2  ;
        PORT
        LAYER M3 ;
        RECT  28.870 249.580 29.600 250.000 ;
        LAYER M2 ;
        RECT  28.870 249.580 29.600 250.000 ;
        END
    END CIN
    PIN OEN
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 80.634  LAYER M2  ;
        ANTENNAPARTIALMETALSIDEAREA 67.374  LAYER M1  ;
        ANTENNAPARTIALMETALSIDEAREA 41.679  LAYER M3  ;
        ANTENNADIFFAREA 0.250  LAYER M3  ;
        ANTENNAPARTIALCUTAREA 0.203  LAYER V2  ;
        ANTENNAPARTIALCUTAREA 0.135  LAYER V3  ;
        ANTENNAGATEAREA 8.100  LAYER M2  ;
        ANTENNAGATEAREA 9.900  LAYER M3  ;
        PORT
        LAYER M3 ;
        RECT  29.900 249.580 30.630 250.000 ;
        LAYER M2 ;
        RECT  29.900 249.580 30.630 250.000 ;
        END
    END OEN
    PIN I
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 67.374  LAYER M1  ;
        ANTENNAPARTIALMETALSIDEAREA 80.804  LAYER M2  ;
        ANTENNAPARTIALMETALSIDEAREA 41.096  LAYER M3  ;
        ANTENNADIFFAREA 0.250  LAYER M3  ;
        ANTENNAPARTIALCUTAREA 0.270  LAYER V2  ;
        ANTENNAPARTIALCUTAREA 0.135  LAYER V3  ;
        ANTENNAGATEAREA 18.900  LAYER M2  ;
        ANTENNAGATEAREA 20.700  LAYER M3  ;
        PORT
        LAYER M3 ;
        RECT  27.840 249.580 28.570 250.000 ;
        LAYER M2 ;
        RECT  27.840 249.580 28.570 250.000 ;
        END
    END I
    PIN VDDO
        DIRECTION INOUT ;
        USE power ;
        PORT
        LAYER M3 ;
        RECT  64.200 192.330 65.000 200.640 ;
        RECT  0.000 201.660 65.000 221.520 ;
        RECT  0.000 222.720 65.000 246.820 ;
        RECT  0.000 192.330 0.800 200.640 ;
        LAYER M2 ;
        RECT  0.000 186.470 65.000 195.650 ;
        LAYER TOP_M ;
        RECT  0.000 195.170 65.000 200.640 ;
        RECT  0.000 201.660 65.000 221.520 ;
        RECT  0.000 222.720 65.000 246.820 ;
        END
    END VDDO
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        PORT
        LAYER M3 ;
        RECT  64.200 163.510 65.000 190.890 ;
        RECT  0.000 163.510 0.800 190.890 ;
        LAYER M2 ;
        RECT  0.000 172.080 65.000 183.060 ;
        LAYER TOP_M ;
        RECT  0.000 163.500 65.000 194.560 ;
        END
    END VDD
    PIN VSSO
        DIRECTION INOUT ;
        USE ground ;
        PORT
        LAYER M3 ;
        RECT  0.000 92.060 65.000 123.250 ;
        RECT  64.200 149.940 65.000 162.610 ;
        RECT  0.000 149.940 0.800 162.610 ;
        LAYER M2 ;
        RECT  0.000 147.040 65.000 154.520 ;
        LAYER TOP_M ;
        RECT  0.000 92.060 65.000 123.250 ;
        RECT  0.000 155.410 65.000 162.610 ;
        END
    END VSSO
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        PORT
        LAYER M3 ;
        RECT  64.200 130.690 65.000 148.880 ;
        RECT  0.000 130.690 0.800 148.880 ;
        LAYER M2 ;
        RECT  0.000 136.310 65.000 146.340 ;
        LAYER TOP_M ;
        RECT  0.000 123.850 65.000 154.560 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  2.000 0.000 63.000 250.000 ;
        RECT  0.000 88.990 65.000 130.360 ;
        RECT  0.000 136.510 65.000 157.550 ;
        RECT  0.315 158.150 64.700 158.460 ;
        RECT  0.300 158.930 64.700 159.230 ;
        RECT  0.300 159.530 64.700 159.830 ;
        RECT  0.300 160.130 64.700 160.430 ;
        RECT  0.300 160.730 64.700 161.030 ;
        RECT  0.300 161.330 64.700 161.630 ;
        RECT  0.300 161.910 64.700 162.190 ;
        RECT  0.300 162.490 64.700 162.770 ;
        RECT  0.300 163.070 64.700 163.350 ;
        RECT  0.300 163.650 64.700 163.950 ;
        RECT  0.300 164.250 64.700 164.550 ;
        RECT  0.300 164.850 64.700 165.150 ;
        RECT  0.300 165.450 64.700 165.750 ;
        RECT  0.300 166.050 64.700 166.350 ;
        RECT  0.300 166.650 64.700 166.960 ;
        RECT  0.300 167.260 64.700 167.560 ;
        RECT  0.300 167.860 64.700 168.160 ;
        RECT  0.000 169.150 65.000 197.240 ;
        RECT  0.600 0.600 64.400 250.000 ;
        RECT  0.000 198.470 65.000 250.000 ;
        LAYER M2 ;
        RECT  1.840 196.420 2.120 249.400 ;
        RECT  63.180 196.430 63.670 249.400 ;
        RECT  0.600 196.440 64.400 245.485 ;
        RECT  26.530 196.440 64.400 248.790 ;
        RECT  0.600 196.440 22.950 249.400 ;
        RECT  26.530 196.440 27.050 249.400 ;
        RECT  31.420 196.440 64.400 249.400 ;
        RECT  19.440 183.720 52.225 185.680 ;
        RECT  0.600 183.850 64.400 185.680 ;
        RECT  46.230 183.720 51.730 185.870 ;
        RECT  55.235 183.850 56.645 185.900 ;
        RECT  4.480 154.920 7.530 171.290 ;
        RECT  8.170 155.125 8.490 171.290 ;
        RECT  22.160 155.160 22.510 171.290 ;
        RECT  22.810 155.140 23.130 171.290 ;
        RECT  31.960 155.120 35.830 171.290 ;
        RECT  49.195 155.130 51.435 171.290 ;
        RECT  52.375 155.300 52.685 171.290 ;
        RECT  53.655 155.035 53.935 171.290 ;
        RECT  56.365 155.280 56.645 171.315 ;
        RECT  57.120 155.300 57.400 171.315 ;
        RECT  57.835 155.130 58.115 171.315 ;
        RECT  0.600 155.310 64.400 171.290 ;
        RECT  56.240 155.310 61.880 171.315 ;
        RECT  53.895 155.310 55.870 171.370 ;
        RECT  3.170 155.310 3.450 171.380 ;
        RECT  34.655 155.310 38.715 171.480 ;
        RECT  39.605 155.310 42.020 171.480 ;
        RECT  2.000 0.000 63.000 60.210 ;
        RECT  0.600 0.600 64.400 60.210 ;
        RECT  0.600 0.600 1.210 135.520 ;
        RECT  0.600 91.020 64.400 135.520 ;
        RECT  4.080 91.020 60.940 135.690 ;
        RECT  62.580 91.020 62.995 135.710 ;
        LAYER M3 ;
        RECT  0.600 247.660 23.220 248.740 ;
        RECT  0.600 247.660 22.900 249.400 ;
        RECT  26.260 247.660 64.400 248.740 ;
        RECT  26.580 247.660 27.000 249.400 ;
        RECT  31.470 247.660 64.400 249.400 ;
        RECT  0.600 124.090 64.400 129.850 ;
        RECT  1.640 124.090 63.600 135.790 ;
        RECT  1.810 124.090 2.830 154.520 ;
        RECT  3.510 124.090 63.600 171.560 ;
        RECT  4.040 123.970 60.900 171.560 ;
        RECT  1.640 155.040 63.600 171.560 ;
        RECT  1.640 183.580 63.600 185.950 ;
        RECT  5.515 124.090 63.600 200.820 ;
        RECT  1.640 196.170 63.600 200.820 ;
        RECT  56.300 123.970 56.580 201.060 ;
        RECT  0.600 0.600 64.400 60.480 ;
        RECT  2.000 0.000 63.000 88.700 ;
        RECT  0.600 0.600 1.480 91.220 ;
        RECT  0.600 90.750 64.400 91.220 ;
        LAYER TOP_M ;
        RECT  0.600 247.690 64.400 248.850 ;
        RECT  0.600 247.690 23.010 249.400 ;
        RECT  26.470 247.690 27.110 249.400 ;
        RECT  31.360 247.690 64.400 249.400 ;
        RECT  2.000 0.000 63.000 91.190 ;
        RECT  0.600 0.600 64.400 91.190 ;
    END
END pt3b03d

MACRO pt3b03
    CLASS PAD ;
    FOREIGN pt3b03 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 65.000 BY 250.000 ;
    SYMMETRY X Y R90 ;
    SITE IOSite_c ;
    PIN PAD
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 55.440  LAYER TOP_M  ;
        ANTENNAPARTIALMETALSIDEAREA 287.938  LAYER M3  ;
        ANTENNAPARTIALMETALSIDEAREA 480.740  LAYER M2  ;
        ANTENNADIFFAREA 2657.280  LAYER TOP_M  ;
        ANTENNADIFFAREA 2657.280  LAYER M3  ;
        ANTENNADIFFAREA 1209.600  LAYER M2  ;
        ANTENNAPARTIALCUTAREA 632.318  LAYER TOP_V  ;
        ANTENNAPARTIALCUTAREA 349.898  LAYER V3  ;
        ANTENNAPARTIALCUTAREA 255.798  LAYER V2  ;
        PORT
        LAYER M3 ;
        RECT  23.740 249.580 25.740 250.000 ;
        LAYER M2 ;
        RECT  2.000 61.000 63.000 90.230 ;
        RECT  23.740 246.275 25.740 250.000 ;
        END
    END PAD
    PIN CIN
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 32.277  LAYER M3  ;
        ANTENNAPARTIALMETALSIDEAREA 96.916  LAYER M2  ;
        ANTENNAPARTIALMETALSIDEAREA 67.374  LAYER M1  ;
        ANTENNADIFFAREA 20.600  LAYER M3  ;
        ANTENNAPARTIALCUTAREA 0.135  LAYER V3  ;
        ANTENNAPARTIALCUTAREA 0.203  LAYER V2  ;
        PORT
        LAYER M3 ;
        RECT  28.870 249.580 29.600 250.000 ;
        LAYER M2 ;
        RECT  28.870 249.580 29.600 250.000 ;
        END
    END CIN
    PIN OEN
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 80.634  LAYER M2  ;
        ANTENNAPARTIALMETALSIDEAREA 67.374  LAYER M1  ;
        ANTENNAPARTIALMETALSIDEAREA 41.679  LAYER M3  ;
        ANTENNADIFFAREA 0.250  LAYER M3  ;
        ANTENNAPARTIALCUTAREA 0.203  LAYER V2  ;
        ANTENNAPARTIALCUTAREA 0.135  LAYER V3  ;
        ANTENNAGATEAREA 8.100  LAYER M2  ;
        ANTENNAGATEAREA 9.900  LAYER M3  ;
        PORT
        LAYER M3 ;
        RECT  29.900 249.580 30.630 250.000 ;
        LAYER M2 ;
        RECT  29.900 249.580 30.630 250.000 ;
        END
    END OEN
    PIN I
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 67.374  LAYER M1  ;
        ANTENNAPARTIALMETALSIDEAREA 80.804  LAYER M2  ;
        ANTENNAPARTIALMETALSIDEAREA 41.096  LAYER M3  ;
        ANTENNADIFFAREA 0.250  LAYER M3  ;
        ANTENNAPARTIALCUTAREA 0.270  LAYER V2  ;
        ANTENNAPARTIALCUTAREA 0.135  LAYER V3  ;
        ANTENNAGATEAREA 18.900  LAYER M2  ;
        ANTENNAGATEAREA 20.700  LAYER M3  ;
        PORT
        LAYER M3 ;
        RECT  27.840 249.580 28.570 250.000 ;
        LAYER M2 ;
        RECT  27.840 249.580 28.570 250.000 ;
        END
    END I
    PIN VDDO
        DIRECTION INOUT ;
        USE power ;
        PORT
        LAYER M3 ;
        RECT  64.200 192.330 65.000 200.640 ;
        RECT  0.000 201.660 65.000 221.520 ;
        RECT  0.000 222.720 65.000 246.820 ;
        RECT  0.000 192.330 0.800 200.640 ;
        LAYER M2 ;
        RECT  0.000 186.470 65.000 195.650 ;
        LAYER TOP_M ;
        RECT  0.000 195.170 65.000 200.640 ;
        RECT  0.000 201.660 65.000 221.520 ;
        RECT  0.000 222.720 65.000 246.820 ;
        END
    END VDDO
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        PORT
        LAYER M3 ;
        RECT  64.200 163.510 65.000 190.890 ;
        RECT  0.000 163.510 0.800 190.890 ;
        LAYER M2 ;
        RECT  0.000 172.080 65.000 183.060 ;
        LAYER TOP_M ;
        RECT  0.000 163.500 65.000 194.560 ;
        END
    END VDD
    PIN VSSO
        DIRECTION INOUT ;
        USE ground ;
        PORT
        LAYER M3 ;
        RECT  0.000 92.060 65.000 123.250 ;
        RECT  64.200 149.940 65.000 162.610 ;
        RECT  0.000 149.940 0.800 162.610 ;
        LAYER M2 ;
        RECT  0.000 147.040 65.000 154.520 ;
        LAYER TOP_M ;
        RECT  0.000 92.060 65.000 123.250 ;
        RECT  0.000 155.410 65.000 162.610 ;
        END
    END VSSO
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        PORT
        LAYER M3 ;
        RECT  64.200 130.690 65.000 148.880 ;
        RECT  0.000 130.690 0.800 148.880 ;
        LAYER M2 ;
        RECT  0.000 136.310 65.000 146.340 ;
        LAYER TOP_M ;
        RECT  0.000 123.850 65.000 154.560 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  2.000 0.000 63.000 250.000 ;
        RECT  0.000 88.990 65.000 130.360 ;
        RECT  0.000 136.510 65.000 157.550 ;
        RECT  0.315 158.150 64.700 158.460 ;
        RECT  0.300 158.930 64.700 159.230 ;
        RECT  0.300 159.530 64.700 159.830 ;
        RECT  0.300 160.130 64.700 160.430 ;
        RECT  0.300 160.730 64.700 161.030 ;
        RECT  0.300 161.330 64.700 161.630 ;
        RECT  0.300 161.910 64.700 162.190 ;
        RECT  0.300 162.490 64.700 162.770 ;
        RECT  0.300 163.070 64.700 163.350 ;
        RECT  0.300 163.650 64.700 163.950 ;
        RECT  0.300 164.250 64.700 164.550 ;
        RECT  0.300 164.850 64.700 165.150 ;
        RECT  0.300 165.450 64.700 165.750 ;
        RECT  0.300 166.050 64.700 166.350 ;
        RECT  0.300 166.650 64.700 166.960 ;
        RECT  0.300 167.260 64.700 167.560 ;
        RECT  0.300 167.860 64.700 168.160 ;
        RECT  0.000 169.150 65.000 197.240 ;
        RECT  0.600 0.600 64.400 250.000 ;
        RECT  0.000 198.470 65.000 250.000 ;
        LAYER M2 ;
        RECT  1.840 196.420 2.120 249.400 ;
        RECT  63.180 196.430 63.670 249.400 ;
        RECT  0.600 196.440 64.400 245.485 ;
        RECT  26.530 196.440 64.400 248.790 ;
        RECT  0.600 196.440 22.950 249.400 ;
        RECT  26.530 196.440 27.050 249.400 ;
        RECT  31.420 196.440 64.400 249.400 ;
        RECT  19.440 183.720 52.225 185.680 ;
        RECT  0.600 183.850 64.400 185.680 ;
        RECT  46.230 183.720 51.730 185.870 ;
        RECT  55.235 183.850 56.645 185.900 ;
        RECT  4.480 154.920 7.530 171.290 ;
        RECT  8.170 155.125 8.490 171.290 ;
        RECT  22.160 155.160 22.510 171.290 ;
        RECT  22.810 155.140 23.130 171.290 ;
        RECT  31.960 155.120 35.830 171.290 ;
        RECT  53.655 155.035 53.935 171.290 ;
        RECT  56.365 155.280 56.645 171.315 ;
        RECT  57.120 155.300 57.400 171.315 ;
        RECT  57.835 155.130 58.115 171.315 ;
        RECT  0.600 155.310 64.400 171.290 ;
        RECT  56.240 155.310 61.880 171.315 ;
        RECT  53.895 155.310 55.870 171.370 ;
        RECT  3.170 155.310 3.450 171.380 ;
        RECT  34.655 155.310 38.715 171.480 ;
        RECT  39.605 155.310 42.020 171.480 ;
        RECT  2.000 0.000 63.000 60.210 ;
        RECT  0.600 0.600 64.400 60.210 ;
        RECT  0.600 0.600 1.210 135.520 ;
        RECT  0.600 91.020 64.400 135.520 ;
        RECT  4.080 91.020 60.940 135.690 ;
        RECT  62.580 91.020 62.995 135.710 ;
        LAYER M3 ;
        RECT  0.600 247.660 23.220 248.740 ;
        RECT  0.600 247.660 22.900 249.400 ;
        RECT  26.260 247.660 64.400 248.740 ;
        RECT  26.580 247.660 27.000 249.400 ;
        RECT  31.470 247.660 64.400 249.400 ;
        RECT  0.600 124.090 64.400 129.850 ;
        RECT  1.640 124.090 63.600 135.790 ;
        RECT  1.810 124.090 2.830 154.520 ;
        RECT  3.510 124.090 63.600 171.560 ;
        RECT  4.040 123.970 60.900 171.560 ;
        RECT  1.640 155.040 63.600 171.560 ;
        RECT  1.640 183.580 63.600 185.950 ;
        RECT  5.515 124.090 63.600 200.820 ;
        RECT  1.640 196.170 63.600 200.820 ;
        RECT  56.300 123.970 56.580 201.060 ;
        RECT  0.600 0.600 64.400 60.480 ;
        RECT  2.000 0.000 63.000 88.700 ;
        RECT  0.600 0.600 1.480 91.220 ;
        RECT  0.600 90.750 64.400 91.220 ;
        LAYER TOP_M ;
        RECT  0.600 247.690 64.400 248.850 ;
        RECT  0.600 247.690 23.010 249.400 ;
        RECT  26.470 247.690 27.110 249.400 ;
        RECT  31.360 247.690 64.400 249.400 ;
        RECT  2.000 0.000 63.000 91.190 ;
        RECT  0.600 0.600 64.400 91.190 ;
    END
END pt3b03

MACRO pt3b02u
    CLASS PAD ;
    FOREIGN pt3b02u 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 65.000 BY 250.000 ;
    SYMMETRY X Y R90 ;
    SITE IOSite_c ;
    PIN PAD
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 55.440  LAYER TOP_M  ;
        ANTENNAPARTIALMETALSIDEAREA 287.938  LAYER M3  ;
        ANTENNAPARTIALMETALSIDEAREA 480.740  LAYER M2  ;
        ANTENNADIFFAREA 2657.280  LAYER TOP_M  ;
        ANTENNADIFFAREA 1209.600  LAYER M2  ;
        ANTENNADIFFAREA 2657.280  LAYER M3  ;
        ANTENNAPARTIALCUTAREA 632.318  LAYER TOP_V  ;
        ANTENNAPARTIALCUTAREA 349.898  LAYER V3  ;
        ANTENNAPARTIALCUTAREA 255.798  LAYER V2  ;
        PORT
        LAYER M3 ;
        RECT  23.740 249.580 25.740 250.000 ;
        LAYER M2 ;
        RECT  2.000 61.000 63.000 90.230 ;
        RECT  23.740 246.275 25.740 250.000 ;
        END
    END PAD
    PIN OEN
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 80.634  LAYER M2  ;
        ANTENNAPARTIALMETALSIDEAREA 41.679  LAYER M3  ;
        ANTENNAPARTIALMETALSIDEAREA 67.374  LAYER M1  ;
        ANTENNADIFFAREA 0.250  LAYER M3  ;
        ANTENNAPARTIALCUTAREA 0.203  LAYER V2  ;
        ANTENNAPARTIALCUTAREA 0.135  LAYER V3  ;
        ANTENNAGATEAREA 9.900  LAYER M3  ;
        ANTENNAGATEAREA 8.100  LAYER M2  ;
        PORT
        LAYER M3 ;
        RECT  29.900 249.580 30.630 250.000 ;
        LAYER M2 ;
        RECT  29.900 249.580 30.630 250.000 ;
        END
    END OEN
    PIN CIN
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 32.277  LAYER M3  ;
        ANTENNAPARTIALMETALSIDEAREA 96.916  LAYER M2  ;
        ANTENNAPARTIALMETALSIDEAREA 67.374  LAYER M1  ;
        ANTENNADIFFAREA 20.600  LAYER M3  ;
        ANTENNAPARTIALCUTAREA 0.135  LAYER V3  ;
        ANTENNAPARTIALCUTAREA 0.203  LAYER V2  ;
        PORT
        LAYER M3 ;
        RECT  28.870 249.580 29.600 250.000 ;
        LAYER M2 ;
        RECT  28.870 249.580 29.600 250.000 ;
        END
    END CIN
    PIN I
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 67.374  LAYER M1  ;
        ANTENNAPARTIALMETALSIDEAREA 80.804  LAYER M2  ;
        ANTENNAPARTIALMETALSIDEAREA 41.096  LAYER M3  ;
        ANTENNADIFFAREA 0.250  LAYER M3  ;
        ANTENNAPARTIALCUTAREA 0.270  LAYER V2  ;
        ANTENNAPARTIALCUTAREA 0.135  LAYER V3  ;
        ANTENNAGATEAREA 18.900  LAYER M2  ;
        ANTENNAGATEAREA 20.700  LAYER M3  ;
        PORT
        LAYER M3 ;
        RECT  27.840 249.580 28.570 250.000 ;
        LAYER M2 ;
        RECT  27.840 249.580 28.570 250.000 ;
        END
    END I
    PIN VDDO
        DIRECTION INOUT ;
        USE power ;
        PORT
        LAYER M3 ;
        RECT  64.200 192.330 65.000 200.640 ;
        RECT  0.000 201.660 65.000 221.520 ;
        RECT  0.000 222.720 65.000 246.820 ;
        RECT  0.000 192.330 0.800 200.640 ;
        LAYER M2 ;
        RECT  0.000 186.470 65.000 195.650 ;
        LAYER TOP_M ;
        RECT  0.000 195.170 65.000 200.640 ;
        RECT  0.000 201.660 65.000 221.520 ;
        RECT  0.000 222.720 65.000 246.820 ;
        END
    END VDDO
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        PORT
        LAYER M3 ;
        RECT  64.200 163.510 65.000 190.890 ;
        RECT  0.000 163.510 0.800 190.890 ;
        LAYER M2 ;
        RECT  0.000 172.080 65.000 183.060 ;
        LAYER TOP_M ;
        RECT  0.000 163.500 65.000 194.560 ;
        END
    END VDD
    PIN VSSO
        DIRECTION INOUT ;
        USE ground ;
        PORT
        LAYER M3 ;
        RECT  0.000 92.060 65.000 123.250 ;
        RECT  64.200 149.940 65.000 162.610 ;
        RECT  0.000 149.940 0.800 162.610 ;
        LAYER M2 ;
        RECT  0.000 147.040 65.000 154.520 ;
        LAYER TOP_M ;
        RECT  0.000 92.060 65.000 123.250 ;
        RECT  0.000 155.410 65.000 162.610 ;
        END
    END VSSO
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        PORT
        LAYER M3 ;
        RECT  64.200 130.690 65.000 148.880 ;
        RECT  0.000 130.690 0.800 148.880 ;
        LAYER M2 ;
        RECT  0.000 136.310 65.000 146.340 ;
        LAYER TOP_M ;
        RECT  0.000 123.850 65.000 154.560 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  2.000 0.000 63.000 250.000 ;
        RECT  0.000 88.990 65.000 130.360 ;
        RECT  0.000 136.510 65.000 157.550 ;
        RECT  0.315 158.150 64.700 158.460 ;
        RECT  0.300 158.930 64.700 159.230 ;
        RECT  0.300 159.530 64.700 159.830 ;
        RECT  0.300 160.130 64.700 160.430 ;
        RECT  0.300 160.730 64.700 161.030 ;
        RECT  0.300 161.330 64.700 161.630 ;
        RECT  0.300 161.910 64.700 162.190 ;
        RECT  0.300 162.490 64.700 162.770 ;
        RECT  0.300 163.070 64.700 163.350 ;
        RECT  0.300 163.650 64.700 163.950 ;
        RECT  0.300 164.250 64.700 164.550 ;
        RECT  0.300 164.850 64.700 165.150 ;
        RECT  0.300 165.450 64.700 165.750 ;
        RECT  0.300 166.050 64.700 166.350 ;
        RECT  0.300 166.650 64.700 166.960 ;
        RECT  0.300 167.260 64.700 167.560 ;
        RECT  0.300 167.860 64.700 168.160 ;
        RECT  0.000 169.150 65.000 197.240 ;
        RECT  0.600 0.600 64.400 250.000 ;
        RECT  0.000 198.470 65.000 250.000 ;
        LAYER M2 ;
        RECT  1.840 196.420 2.120 249.400 ;
        RECT  63.180 196.430 63.670 249.400 ;
        RECT  0.600 196.440 64.400 245.485 ;
        RECT  26.530 196.440 64.400 248.790 ;
        RECT  0.600 196.440 22.950 249.400 ;
        RECT  26.530 196.440 27.050 249.400 ;
        RECT  31.420 196.440 64.400 249.400 ;
        RECT  19.440 183.720 52.185 185.680 ;
        RECT  0.600 183.850 64.400 185.680 ;
        RECT  46.230 183.720 51.730 185.870 ;
        RECT  54.855 183.850 56.700 185.950 ;
        RECT  4.895 155.120 7.525 171.290 ;
        RECT  8.170 155.125 8.490 171.290 ;
        RECT  22.160 155.160 22.510 171.290 ;
        RECT  22.810 155.140 23.130 171.290 ;
        RECT  53.655 155.035 53.935 171.290 ;
        RECT  56.365 155.280 56.645 171.315 ;
        RECT  57.120 155.300 57.400 171.315 ;
        RECT  57.835 155.130 58.115 171.315 ;
        RECT  0.600 155.310 64.400 171.290 ;
        RECT  56.240 155.310 61.880 171.315 ;
        RECT  33.625 155.310 34.125 171.365 ;
        RECT  53.895 155.310 55.870 171.370 ;
        RECT  3.220 155.310 3.500 171.380 ;
        RECT  34.655 155.310 38.715 171.480 ;
        RECT  39.605 155.310 42.020 171.480 ;
        RECT  2.000 0.000 63.000 60.210 ;
        RECT  0.600 0.600 64.400 60.210 ;
        RECT  0.600 0.600 1.210 135.520 ;
        RECT  0.600 91.020 64.400 135.520 ;
        RECT  4.080 91.020 60.940 135.690 ;
        RECT  62.580 91.020 62.995 135.710 ;
        LAYER M3 ;
        RECT  0.600 247.660 23.220 248.740 ;
        RECT  0.600 247.660 22.900 249.400 ;
        RECT  26.260 247.660 64.400 248.740 ;
        RECT  26.580 247.660 27.000 249.400 ;
        RECT  31.470 247.660 64.400 249.400 ;
        RECT  0.600 124.090 64.400 129.850 ;
        RECT  1.640 124.090 63.600 135.790 ;
        RECT  1.810 124.090 2.830 154.520 ;
        RECT  3.110 124.090 63.600 171.560 ;
        RECT  4.040 123.970 60.900 171.560 ;
        RECT  1.640 155.040 63.600 171.560 ;
        RECT  1.640 183.580 63.600 185.950 ;
        RECT  5.510 124.090 63.600 200.820 ;
        RECT  1.640 196.170 63.600 200.820 ;
        RECT  56.300 123.970 56.580 201.060 ;
        RECT  0.600 0.600 64.400 60.480 ;
        RECT  2.000 0.000 63.000 88.700 ;
        RECT  0.600 0.600 1.480 91.220 ;
        RECT  0.600 90.750 64.400 91.220 ;
        LAYER TOP_M ;
        RECT  0.600 247.690 64.400 248.850 ;
        RECT  0.600 247.690 23.010 249.400 ;
        RECT  26.470 247.690 27.110 249.400 ;
        RECT  31.360 247.690 64.400 249.400 ;
        RECT  2.000 0.000 63.000 91.190 ;
        RECT  0.600 0.600 64.400 91.190 ;
    END
END pt3b02u

MACRO pt3b02d
    CLASS PAD ;
    FOREIGN pt3b02d 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 65.000 BY 250.000 ;
    SYMMETRY X Y R90 ;
    SITE IOSite_c ;
    PIN PAD
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 55.440  LAYER TOP_M  ;
        ANTENNAPARTIALMETALSIDEAREA 287.938  LAYER M3  ;
        ANTENNAPARTIALMETALSIDEAREA 480.740  LAYER M2  ;
        ANTENNADIFFAREA 2657.280  LAYER TOP_M  ;
        ANTENNADIFFAREA 1209.600  LAYER M2  ;
        ANTENNADIFFAREA 2657.280  LAYER M3  ;
        ANTENNAPARTIALCUTAREA 632.318  LAYER TOP_V  ;
        ANTENNAPARTIALCUTAREA 349.898  LAYER V3  ;
        ANTENNAPARTIALCUTAREA 255.798  LAYER V2  ;
        PORT
        LAYER M3 ;
        RECT  23.740 249.580 25.740 250.000 ;
        LAYER M2 ;
        RECT  2.000 61.000 63.000 90.230 ;
        RECT  23.740 246.275 25.740 250.000 ;
        END
    END PAD
    PIN OEN
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 80.634  LAYER M2  ;
        ANTENNAPARTIALMETALSIDEAREA 41.679  LAYER M3  ;
        ANTENNAPARTIALMETALSIDEAREA 67.374  LAYER M1  ;
        ANTENNADIFFAREA 0.250  LAYER M3  ;
        ANTENNAPARTIALCUTAREA 0.203  LAYER V2  ;
        ANTENNAPARTIALCUTAREA 0.135  LAYER V3  ;
        ANTENNAGATEAREA 9.900  LAYER M3  ;
        ANTENNAGATEAREA 8.100  LAYER M2  ;
        PORT
        LAYER M3 ;
        RECT  29.900 249.580 30.630 250.000 ;
        LAYER M2 ;
        RECT  29.900 249.580 30.630 250.000 ;
        END
    END OEN
    PIN CIN
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 32.277  LAYER M3  ;
        ANTENNAPARTIALMETALSIDEAREA 96.916  LAYER M2  ;
        ANTENNAPARTIALMETALSIDEAREA 67.374  LAYER M1  ;
        ANTENNADIFFAREA 20.600  LAYER M3  ;
        ANTENNAPARTIALCUTAREA 0.135  LAYER V3  ;
        ANTENNAPARTIALCUTAREA 0.203  LAYER V2  ;
        PORT
        LAYER M3 ;
        RECT  28.870 249.580 29.600 250.000 ;
        LAYER M2 ;
        RECT  28.870 249.580 29.600 250.000 ;
        END
    END CIN
    PIN I
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 67.374  LAYER M1  ;
        ANTENNAPARTIALMETALSIDEAREA 80.804  LAYER M2  ;
        ANTENNAPARTIALMETALSIDEAREA 41.096  LAYER M3  ;
        ANTENNADIFFAREA 0.250  LAYER M3  ;
        ANTENNAPARTIALCUTAREA 0.270  LAYER V2  ;
        ANTENNAPARTIALCUTAREA 0.135  LAYER V3  ;
        ANTENNAGATEAREA 18.900  LAYER M2  ;
        ANTENNAGATEAREA 20.700  LAYER M3  ;
        PORT
        LAYER M3 ;
        RECT  27.840 249.580 28.570 250.000 ;
        LAYER M2 ;
        RECT  27.840 249.580 28.570 250.000 ;
        END
    END I
    PIN VDDO
        DIRECTION INOUT ;
        USE power ;
        PORT
        LAYER M3 ;
        RECT  64.200 192.330 65.000 200.640 ;
        RECT  0.000 201.660 65.000 221.520 ;
        RECT  0.000 222.720 65.000 246.820 ;
        RECT  0.000 192.330 0.800 200.640 ;
        LAYER M2 ;
        RECT  0.000 186.470 65.000 195.650 ;
        LAYER TOP_M ;
        RECT  0.000 195.170 65.000 200.640 ;
        RECT  0.000 201.660 65.000 221.520 ;
        RECT  0.000 222.720 65.000 246.820 ;
        END
    END VDDO
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        PORT
        LAYER M3 ;
        RECT  64.200 163.510 65.000 190.890 ;
        RECT  0.000 163.510 0.800 190.890 ;
        LAYER M2 ;
        RECT  0.000 172.080 65.000 183.060 ;
        LAYER TOP_M ;
        RECT  0.000 163.500 65.000 194.560 ;
        END
    END VDD
    PIN VSSO
        DIRECTION INOUT ;
        USE ground ;
        PORT
        LAYER M3 ;
        RECT  0.000 92.060 65.000 123.250 ;
        RECT  64.200 149.940 65.000 162.610 ;
        RECT  0.000 149.940 0.800 162.610 ;
        LAYER M2 ;
        RECT  0.000 147.040 65.000 154.520 ;
        LAYER TOP_M ;
        RECT  0.000 92.060 65.000 123.250 ;
        RECT  0.000 155.410 65.000 162.610 ;
        END
    END VSSO
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        PORT
        LAYER M3 ;
        RECT  64.200 130.690 65.000 148.880 ;
        RECT  0.000 130.690 0.800 148.880 ;
        LAYER M2 ;
        RECT  0.000 136.310 65.000 146.340 ;
        LAYER TOP_M ;
        RECT  0.000 123.850 65.000 154.560 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  2.000 0.000 63.000 250.000 ;
        RECT  0.000 88.990 65.000 130.360 ;
        RECT  0.000 136.510 65.000 157.550 ;
        RECT  0.315 158.150 64.700 158.460 ;
        RECT  0.300 158.930 64.700 159.230 ;
        RECT  0.300 159.530 64.700 159.830 ;
        RECT  0.300 160.130 64.700 160.430 ;
        RECT  0.300 160.730 64.700 161.030 ;
        RECT  0.300 161.330 64.700 161.630 ;
        RECT  0.300 161.910 64.700 162.190 ;
        RECT  0.300 162.490 64.700 162.770 ;
        RECT  0.300 163.070 64.700 163.350 ;
        RECT  0.300 163.650 64.700 163.950 ;
        RECT  0.300 164.250 64.700 164.550 ;
        RECT  0.300 164.850 64.700 165.150 ;
        RECT  0.300 165.450 64.700 165.750 ;
        RECT  0.300 166.050 64.700 166.350 ;
        RECT  0.300 166.650 64.700 166.960 ;
        RECT  0.300 167.260 64.700 167.560 ;
        RECT  0.300 167.860 64.700 168.160 ;
        RECT  0.000 169.150 65.000 197.240 ;
        RECT  0.600 0.600 64.400 250.000 ;
        RECT  0.000 198.470 65.000 250.000 ;
        LAYER M2 ;
        RECT  1.840 196.420 2.120 249.400 ;
        RECT  63.180 196.430 63.670 249.400 ;
        RECT  0.600 196.440 64.400 245.485 ;
        RECT  26.530 196.440 64.400 248.790 ;
        RECT  0.600 196.440 22.950 249.400 ;
        RECT  26.530 196.440 27.050 249.400 ;
        RECT  31.420 196.440 64.400 249.400 ;
        RECT  19.440 183.720 52.185 185.680 ;
        RECT  0.600 183.850 64.400 185.680 ;
        RECT  46.230 183.720 51.730 185.870 ;
        RECT  54.855 183.850 56.700 185.950 ;
        RECT  4.895 155.120 7.525 171.290 ;
        RECT  8.170 155.125 8.490 171.290 ;
        RECT  22.160 155.160 22.510 171.290 ;
        RECT  22.810 155.140 23.130 171.290 ;
        RECT  49.620 155.125 51.860 171.290 ;
        RECT  52.800 155.295 53.110 171.290 ;
        RECT  53.655 155.035 53.935 171.290 ;
        RECT  56.365 155.280 56.645 171.315 ;
        RECT  57.120 155.300 57.400 171.315 ;
        RECT  57.835 155.130 58.115 171.315 ;
        RECT  0.600 155.310 64.400 171.290 ;
        RECT  56.240 155.310 61.880 171.315 ;
        RECT  53.895 155.310 55.870 171.370 ;
        RECT  3.220 155.310 3.500 171.380 ;
        RECT  34.655 155.310 38.715 171.480 ;
        RECT  39.605 155.310 42.020 171.480 ;
        RECT  2.000 0.000 63.000 60.210 ;
        RECT  0.600 0.600 64.400 60.210 ;
        RECT  0.600 0.600 1.210 135.520 ;
        RECT  0.600 91.020 64.400 135.520 ;
        RECT  4.080 91.020 60.940 135.690 ;
        RECT  62.580 91.020 62.995 135.710 ;
        LAYER M3 ;
        RECT  0.600 247.660 23.220 248.740 ;
        RECT  0.600 247.660 22.900 249.400 ;
        RECT  26.260 247.660 64.400 248.740 ;
        RECT  26.580 247.660 27.000 249.400 ;
        RECT  31.470 247.660 64.400 249.400 ;
        RECT  0.600 124.090 64.400 129.850 ;
        RECT  1.640 124.090 63.600 135.790 ;
        RECT  1.810 124.090 2.830 154.520 ;
        RECT  3.110 124.090 63.600 171.560 ;
        RECT  4.040 123.970 60.900 171.560 ;
        RECT  1.640 155.040 63.600 171.560 ;
        RECT  1.640 183.580 63.600 185.950 ;
        RECT  5.510 124.090 63.600 200.820 ;
        RECT  1.640 196.170 63.600 200.820 ;
        RECT  56.300 123.970 56.580 201.060 ;
        RECT  0.600 0.600 64.400 60.480 ;
        RECT  2.000 0.000 63.000 88.700 ;
        RECT  0.600 0.600 1.480 91.220 ;
        RECT  0.600 90.750 64.400 91.220 ;
        LAYER TOP_M ;
        RECT  0.600 247.690 64.400 248.850 ;
        RECT  0.600 247.690 23.010 249.400 ;
        RECT  26.470 247.690 27.110 249.400 ;
        RECT  31.360 247.690 64.400 249.400 ;
        RECT  2.000 0.000 63.000 91.190 ;
        RECT  0.600 0.600 64.400 91.190 ;
    END
END pt3b02d

MACRO pt3b02
    CLASS PAD ;
    FOREIGN pt3b02 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 65.000 BY 250.000 ;
    SYMMETRY X Y R90 ;
    SITE IOSite_c ;
    PIN PAD
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 55.440  LAYER TOP_M  ;
        ANTENNAPARTIALMETALSIDEAREA 287.938  LAYER M3  ;
        ANTENNAPARTIALMETALSIDEAREA 480.740  LAYER M2  ;
        ANTENNADIFFAREA 2657.280  LAYER TOP_M  ;
        ANTENNADIFFAREA 1209.600  LAYER M2  ;
        ANTENNADIFFAREA 2657.280  LAYER M3  ;
        ANTENNAPARTIALCUTAREA 632.318  LAYER TOP_V  ;
        ANTENNAPARTIALCUTAREA 349.898  LAYER V3  ;
        ANTENNAPARTIALCUTAREA 255.798  LAYER V2  ;
        PORT
        LAYER M3 ;
        RECT  23.740 249.580 25.740 250.000 ;
        LAYER M2 ;
        RECT  2.000 61.000 63.000 90.230 ;
        RECT  23.740 246.275 25.740 250.000 ;
        END
    END PAD
    PIN OEN
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 80.634  LAYER M2  ;
        ANTENNAPARTIALMETALSIDEAREA 41.679  LAYER M3  ;
        ANTENNAPARTIALMETALSIDEAREA 67.374  LAYER M1  ;
        ANTENNADIFFAREA 0.250  LAYER M3  ;
        ANTENNAPARTIALCUTAREA 0.203  LAYER V2  ;
        ANTENNAPARTIALCUTAREA 0.135  LAYER V3  ;
        ANTENNAGATEAREA 9.900  LAYER M3  ;
        ANTENNAGATEAREA 8.100  LAYER M2  ;
        PORT
        LAYER M3 ;
        RECT  29.900 249.580 30.630 250.000 ;
        LAYER M2 ;
        RECT  29.900 249.580 30.630 250.000 ;
        END
    END OEN
    PIN CIN
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 32.277  LAYER M3  ;
        ANTENNAPARTIALMETALSIDEAREA 96.916  LAYER M2  ;
        ANTENNAPARTIALMETALSIDEAREA 67.374  LAYER M1  ;
        ANTENNADIFFAREA 20.600  LAYER M3  ;
        ANTENNAPARTIALCUTAREA 0.135  LAYER V3  ;
        ANTENNAPARTIALCUTAREA 0.203  LAYER V2  ;
        PORT
        LAYER M3 ;
        RECT  28.870 249.580 29.600 250.000 ;
        LAYER M2 ;
        RECT  28.870 249.580 29.600 250.000 ;
        END
    END CIN
    PIN I
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 67.374  LAYER M1  ;
        ANTENNAPARTIALMETALSIDEAREA 80.804  LAYER M2  ;
        ANTENNAPARTIALMETALSIDEAREA 41.096  LAYER M3  ;
        ANTENNADIFFAREA 0.250  LAYER M3  ;
        ANTENNAPARTIALCUTAREA 0.270  LAYER V2  ;
        ANTENNAPARTIALCUTAREA 0.135  LAYER V3  ;
        ANTENNAGATEAREA 18.900  LAYER M2  ;
        ANTENNAGATEAREA 20.700  LAYER M3  ;
        PORT
        LAYER M3 ;
        RECT  27.840 249.580 28.570 250.000 ;
        LAYER M2 ;
        RECT  27.840 249.580 28.570 250.000 ;
        END
    END I
    PIN VDDO
        DIRECTION INOUT ;
        USE power ;
        PORT
        LAYER M3 ;
        RECT  64.200 192.330 65.000 200.640 ;
        RECT  0.000 201.660 65.000 221.520 ;
        RECT  0.000 222.720 65.000 246.820 ;
        RECT  0.000 192.330 0.800 200.640 ;
        LAYER M2 ;
        RECT  0.000 186.470 65.000 195.650 ;
        LAYER TOP_M ;
        RECT  0.000 195.170 65.000 200.640 ;
        RECT  0.000 201.660 65.000 221.520 ;
        RECT  0.000 222.720 65.000 246.820 ;
        END
    END VDDO
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        PORT
        LAYER M3 ;
        RECT  64.200 163.510 65.000 190.890 ;
        RECT  0.000 163.510 0.800 190.890 ;
        LAYER M2 ;
        RECT  0.000 172.080 65.000 183.060 ;
        LAYER TOP_M ;
        RECT  0.000 163.500 65.000 194.560 ;
        END
    END VDD
    PIN VSSO
        DIRECTION INOUT ;
        USE ground ;
        PORT
        LAYER M3 ;
        RECT  0.000 92.060 65.000 123.250 ;
        RECT  64.200 149.940 65.000 162.610 ;
        RECT  0.000 149.940 0.800 162.610 ;
        LAYER M2 ;
        RECT  0.000 147.040 65.000 154.520 ;
        LAYER TOP_M ;
        RECT  0.000 92.060 65.000 123.250 ;
        RECT  0.000 155.410 65.000 162.610 ;
        END
    END VSSO
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        PORT
        LAYER M3 ;
        RECT  64.200 130.690 65.000 148.880 ;
        RECT  0.000 130.690 0.800 148.880 ;
        LAYER M2 ;
        RECT  0.000 136.310 65.000 146.340 ;
        LAYER TOP_M ;
        RECT  0.000 123.850 65.000 154.560 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  2.000 0.000 63.000 250.000 ;
        RECT  0.000 88.990 65.000 130.360 ;
        RECT  0.000 136.510 65.000 157.550 ;
        RECT  0.315 158.150 64.700 158.460 ;
        RECT  0.300 158.930 64.700 159.230 ;
        RECT  0.300 159.530 64.700 159.830 ;
        RECT  0.300 160.130 64.700 160.430 ;
        RECT  0.300 160.730 64.700 161.030 ;
        RECT  0.300 161.330 64.700 161.630 ;
        RECT  0.300 161.910 64.700 162.190 ;
        RECT  0.300 162.490 64.700 162.770 ;
        RECT  0.300 163.070 64.700 163.350 ;
        RECT  0.300 163.650 64.700 163.950 ;
        RECT  0.300 164.250 64.700 164.550 ;
        RECT  0.300 164.850 64.700 165.150 ;
        RECT  0.300 165.450 64.700 165.750 ;
        RECT  0.300 166.050 64.700 166.350 ;
        RECT  0.300 166.650 64.700 166.960 ;
        RECT  0.300 167.260 64.700 167.560 ;
        RECT  0.300 167.860 64.700 168.160 ;
        RECT  0.000 169.150 65.000 197.240 ;
        RECT  0.600 0.600 64.400 250.000 ;
        RECT  0.000 198.470 65.000 250.000 ;
        LAYER M2 ;
        RECT  1.840 196.420 2.120 249.400 ;
        RECT  63.180 196.430 63.670 249.400 ;
        RECT  0.600 196.440 64.400 245.485 ;
        RECT  26.530 196.440 64.400 248.790 ;
        RECT  0.600 196.440 22.950 249.400 ;
        RECT  26.530 196.440 27.050 249.400 ;
        RECT  31.420 196.440 64.400 249.400 ;
        RECT  19.440 183.720 52.185 185.680 ;
        RECT  0.600 183.850 64.400 185.680 ;
        RECT  46.230 183.720 51.730 185.870 ;
        RECT  54.855 183.850 56.700 185.950 ;
        RECT  4.895 155.120 7.525 171.290 ;
        RECT  8.170 155.125 8.490 171.290 ;
        RECT  22.160 155.160 22.510 171.290 ;
        RECT  22.810 155.140 23.130 171.290 ;
        RECT  53.655 155.035 53.935 171.290 ;
        RECT  56.365 155.280 56.645 171.315 ;
        RECT  57.120 155.300 57.400 171.315 ;
        RECT  57.835 155.130 58.115 171.315 ;
        RECT  0.600 155.310 64.400 171.290 ;
        RECT  56.240 155.310 61.880 171.315 ;
        RECT  53.895 155.310 55.870 171.370 ;
        RECT  3.220 155.310 3.500 171.380 ;
        RECT  34.655 155.310 38.715 171.480 ;
        RECT  39.605 155.310 42.020 171.480 ;
        RECT  2.000 0.000 63.000 60.210 ;
        RECT  0.600 0.600 64.400 60.210 ;
        RECT  0.600 0.600 1.210 135.520 ;
        RECT  0.600 91.020 64.400 135.520 ;
        RECT  4.080 91.020 60.940 135.690 ;
        RECT  62.580 91.020 62.995 135.710 ;
        LAYER M3 ;
        RECT  0.600 247.660 23.220 248.740 ;
        RECT  0.600 247.660 22.900 249.400 ;
        RECT  26.260 247.660 64.400 248.740 ;
        RECT  26.580 247.660 27.000 249.400 ;
        RECT  31.470 247.660 64.400 249.400 ;
        RECT  0.600 124.090 64.400 129.850 ;
        RECT  1.640 124.090 63.600 135.790 ;
        RECT  1.810 124.090 2.830 154.520 ;
        RECT  3.110 124.090 63.600 171.560 ;
        RECT  4.040 123.970 60.900 171.560 ;
        RECT  1.640 155.040 63.600 171.560 ;
        RECT  1.640 183.580 63.600 185.950 ;
        RECT  5.510 124.090 63.600 200.820 ;
        RECT  1.640 196.170 63.600 200.820 ;
        RECT  56.300 123.970 56.580 201.060 ;
        RECT  0.600 0.600 64.400 60.480 ;
        RECT  2.000 0.000 63.000 88.700 ;
        RECT  0.600 0.600 1.480 91.220 ;
        RECT  0.600 90.750 64.400 91.220 ;
        LAYER TOP_M ;
        RECT  0.600 247.690 64.400 248.850 ;
        RECT  0.600 247.690 23.010 249.400 ;
        RECT  26.470 247.690 27.110 249.400 ;
        RECT  31.360 247.690 64.400 249.400 ;
        RECT  2.000 0.000 63.000 91.190 ;
        RECT  0.600 0.600 64.400 91.190 ;
    END
END pt3b02

MACRO pt3b01u
    CLASS PAD ;
    FOREIGN pt3b01u 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 65.000 BY 250.000 ;
    SYMMETRY X Y R90 ;
    SITE IOSite_c ;
    PIN PAD
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 55.440  LAYER TOP_M  ;
        ANTENNAPARTIALMETALSIDEAREA 287.938  LAYER M3  ;
        ANTENNAPARTIALMETALSIDEAREA 480.740  LAYER M2  ;
        ANTENNADIFFAREA 2657.280  LAYER TOP_M  ;
        ANTENNADIFFAREA 2657.280  LAYER M3  ;
        ANTENNADIFFAREA 1209.600  LAYER M2  ;
        ANTENNAPARTIALCUTAREA 632.318  LAYER TOP_V  ;
        ANTENNAPARTIALCUTAREA 349.898  LAYER V3  ;
        ANTENNAPARTIALCUTAREA 255.798  LAYER V2  ;
        PORT
        LAYER M3 ;
        RECT  23.740 249.580 25.740 250.000 ;
        LAYER M2 ;
        RECT  2.000 61.000 63.000 90.230 ;
        RECT  23.740 246.275 25.740 250.000 ;
        END
    END PAD
    PIN OEN
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 67.374  LAYER M1  ;
        ANTENNAPARTIALMETALSIDEAREA 80.634  LAYER M2  ;
        ANTENNAPARTIALMETALSIDEAREA 41.679  LAYER M3  ;
        ANTENNADIFFAREA 0.250  LAYER M3  ;
        ANTENNAPARTIALCUTAREA 0.203  LAYER V2  ;
        ANTENNAPARTIALCUTAREA 0.135  LAYER V3  ;
        ANTENNAGATEAREA 8.100  LAYER M2  ;
        ANTENNAGATEAREA 9.900  LAYER M3  ;
        PORT
        LAYER M3 ;
        RECT  29.900 249.580 30.630 250.000 ;
        LAYER M2 ;
        RECT  29.900 249.580 30.630 250.000 ;
        END
    END OEN
    PIN CIN
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 32.277  LAYER M3  ;
        ANTENNAPARTIALMETALSIDEAREA 96.916  LAYER M2  ;
        ANTENNAPARTIALMETALSIDEAREA 67.374  LAYER M1  ;
        ANTENNADIFFAREA 20.600  LAYER M3  ;
        ANTENNAPARTIALCUTAREA 0.135  LAYER V3  ;
        ANTENNAPARTIALCUTAREA 0.203  LAYER V2  ;
        PORT
        LAYER M3 ;
        RECT  28.870 249.580 29.600 250.000 ;
        LAYER M2 ;
        RECT  28.870 249.580 29.600 250.000 ;
        END
    END CIN
    PIN I
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 80.804  LAYER M2  ;
        ANTENNAPARTIALMETALSIDEAREA 67.374  LAYER M1  ;
        ANTENNAPARTIALMETALSIDEAREA 41.096  LAYER M3  ;
        ANTENNADIFFAREA 0.250  LAYER M3  ;
        ANTENNAPARTIALCUTAREA 0.203  LAYER V2  ;
        ANTENNAPARTIALCUTAREA 0.135  LAYER V3  ;
        ANTENNAGATEAREA 8.100  LAYER M2  ;
        ANTENNAGATEAREA 9.900  LAYER M3  ;
        PORT
        LAYER M3 ;
        RECT  27.840 249.580 28.570 250.000 ;
        LAYER M2 ;
        RECT  27.840 249.580 28.570 250.000 ;
        END
    END I
    PIN VDDO
        DIRECTION INOUT ;
        USE power ;
        PORT
        LAYER M3 ;
        RECT  64.200 192.330 65.000 200.640 ;
        RECT  0.000 201.660 65.000 221.520 ;
        RECT  0.000 222.720 65.000 246.820 ;
        RECT  0.000 192.330 0.800 200.640 ;
        LAYER M2 ;
        RECT  0.000 186.470 65.000 195.650 ;
        LAYER TOP_M ;
        RECT  0.000 195.170 65.000 200.640 ;
        RECT  0.000 201.660 65.000 221.520 ;
        RECT  0.000 222.720 65.000 246.820 ;
        END
    END VDDO
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        PORT
        LAYER M3 ;
        RECT  64.200 163.510 65.000 190.890 ;
        RECT  0.000 163.510 0.800 190.890 ;
        LAYER M2 ;
        RECT  0.000 172.080 65.000 183.060 ;
        LAYER TOP_M ;
        RECT  0.000 163.500 65.000 194.560 ;
        END
    END VDD
    PIN VSSO
        DIRECTION INOUT ;
        USE ground ;
        PORT
        LAYER M3 ;
        RECT  0.000 92.060 65.000 123.250 ;
        RECT  64.200 149.940 65.000 162.610 ;
        RECT  0.000 149.940 0.800 162.610 ;
        LAYER M2 ;
        RECT  0.000 147.040 65.000 154.520 ;
        LAYER TOP_M ;
        RECT  0.000 92.060 65.000 123.250 ;
        RECT  0.000 155.410 65.000 162.610 ;
        END
    END VSSO
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        PORT
        LAYER M3 ;
        RECT  64.200 130.690 65.000 148.880 ;
        RECT  0.000 130.690 0.800 148.880 ;
        LAYER M2 ;
        RECT  0.000 136.310 65.000 146.340 ;
        LAYER TOP_M ;
        RECT  0.000 123.850 65.000 154.560 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  2.000 0.000 63.000 250.000 ;
        RECT  0.000 88.990 65.000 130.360 ;
        RECT  0.000 136.510 65.000 157.550 ;
        RECT  0.315 158.150 64.700 158.460 ;
        RECT  0.300 158.930 64.700 159.230 ;
        RECT  0.300 159.530 64.700 159.830 ;
        RECT  0.300 160.130 64.700 160.430 ;
        RECT  0.300 160.730 64.700 161.030 ;
        RECT  0.300 161.330 64.700 161.630 ;
        RECT  0.300 161.910 64.700 162.190 ;
        RECT  0.300 162.490 64.700 162.770 ;
        RECT  0.300 163.070 64.700 163.350 ;
        RECT  0.300 163.650 64.700 163.950 ;
        RECT  0.300 164.250 64.700 164.550 ;
        RECT  0.300 164.850 64.700 165.150 ;
        RECT  0.300 165.450 64.700 165.750 ;
        RECT  0.300 166.050 64.700 166.350 ;
        RECT  0.300 166.650 64.700 166.960 ;
        RECT  0.300 167.260 64.700 167.560 ;
        RECT  0.300 167.860 64.700 168.160 ;
        RECT  0.000 169.150 65.000 197.240 ;
        RECT  0.600 0.600 64.400 250.000 ;
        RECT  0.000 198.470 65.000 250.000 ;
        LAYER M2 ;
        RECT  1.840 196.420 2.120 249.400 ;
        RECT  63.180 196.430 63.670 249.400 ;
        RECT  0.600 196.440 64.400 245.485 ;
        RECT  26.530 196.440 64.400 248.790 ;
        RECT  0.600 196.440 22.950 249.400 ;
        RECT  26.530 196.440 27.050 249.400 ;
        RECT  31.420 196.440 64.400 249.400 ;
        RECT  14.290 183.720 52.380 185.680 ;
        RECT  0.600 183.850 64.400 185.680 ;
        RECT  54.910 183.850 57.160 185.865 ;
        RECT  46.230 183.720 51.730 185.870 ;
        RECT  18.450 155.160 18.800 171.290 ;
        RECT  19.100 155.140 19.420 171.290 ;
        RECT  53.655 155.035 53.935 171.290 ;
        RECT  56.365 155.280 56.645 171.315 ;
        RECT  57.120 155.300 57.400 171.315 ;
        RECT  57.835 155.130 58.115 171.315 ;
        RECT  0.600 155.310 64.400 171.290 ;
        RECT  56.240 155.310 61.880 171.315 ;
        RECT  53.895 155.310 55.870 171.370 ;
        RECT  31.880 155.310 32.380 171.375 ;
        RECT  3.210 155.310 3.490 171.380 ;
        RECT  34.655 155.310 38.715 171.480 ;
        RECT  39.605 155.310 42.020 171.480 ;
        RECT  2.000 0.000 63.000 60.210 ;
        RECT  0.600 0.600 64.400 60.210 ;
        RECT  0.600 0.600 1.210 135.520 ;
        RECT  0.600 91.020 64.400 135.520 ;
        RECT  4.080 91.020 60.940 135.690 ;
        RECT  62.580 91.020 62.995 135.710 ;
        LAYER M3 ;
        RECT  0.600 247.660 23.220 248.740 ;
        RECT  0.600 247.660 22.900 249.400 ;
        RECT  26.260 247.660 64.400 248.740 ;
        RECT  26.580 247.660 27.000 249.400 ;
        RECT  31.470 247.660 64.400 249.400 ;
        RECT  0.600 124.090 64.400 129.850 ;
        RECT  3.990 123.970 60.900 135.790 ;
        RECT  1.640 124.090 63.600 135.790 ;
        RECT  1.810 124.090 2.830 154.520 ;
        RECT  5.155 123.970 60.900 171.560 ;
        RECT  1.640 155.040 63.600 171.560 ;
        RECT  1.640 183.580 63.600 185.950 ;
        RECT  5.490 124.090 63.600 200.820 ;
        RECT  1.640 196.170 63.600 200.820 ;
        RECT  56.300 123.970 56.580 201.060 ;
        RECT  0.600 0.600 64.400 60.480 ;
        RECT  2.000 0.000 63.000 88.700 ;
        RECT  0.600 0.600 1.480 91.220 ;
        RECT  0.600 90.750 64.400 91.220 ;
        LAYER TOP_M ;
        RECT  0.600 247.690 64.400 248.850 ;
        RECT  0.600 247.690 23.010 249.400 ;
        RECT  26.470 247.690 27.110 249.400 ;
        RECT  31.360 247.690 64.400 249.400 ;
        RECT  2.000 0.000 63.000 91.190 ;
        RECT  0.600 0.600 64.400 91.190 ;
    END
END pt3b01u

MACRO pt3b01d
    CLASS PAD ;
    FOREIGN pt3b01d 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 65.000 BY 250.000 ;
    SYMMETRY X Y R90 ;
    SITE IOSite_c ;
    PIN PAD
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 55.440  LAYER TOP_M  ;
        ANTENNAPARTIALMETALSIDEAREA 287.938  LAYER M3  ;
        ANTENNAPARTIALMETALSIDEAREA 480.740  LAYER M2  ;
        ANTENNADIFFAREA 2657.280  LAYER TOP_M  ;
        ANTENNADIFFAREA 2657.280  LAYER M3  ;
        ANTENNADIFFAREA 1209.600  LAYER M2  ;
        ANTENNAPARTIALCUTAREA 632.318  LAYER TOP_V  ;
        ANTENNAPARTIALCUTAREA 349.898  LAYER V3  ;
        ANTENNAPARTIALCUTAREA 255.798  LAYER V2  ;
        PORT
        LAYER M3 ;
        RECT  23.740 249.580 25.740 250.000 ;
        LAYER M2 ;
        RECT  2.000 61.000 63.000 90.230 ;
        RECT  23.740 246.275 25.740 250.000 ;
        END
    END PAD
    PIN OEN
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 67.374  LAYER M1  ;
        ANTENNAPARTIALMETALSIDEAREA 80.634  LAYER M2  ;
        ANTENNAPARTIALMETALSIDEAREA 41.679  LAYER M3  ;
        ANTENNADIFFAREA 0.250  LAYER M3  ;
        ANTENNAPARTIALCUTAREA 0.203  LAYER V2  ;
        ANTENNAPARTIALCUTAREA 0.135  LAYER V3  ;
        ANTENNAGATEAREA 8.100  LAYER M2  ;
        ANTENNAGATEAREA 9.900  LAYER M3  ;
        PORT
        LAYER M3 ;
        RECT  29.900 249.580 30.630 250.000 ;
        LAYER M2 ;
        RECT  29.900 249.580 30.630 250.000 ;
        END
    END OEN
    PIN CIN
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 32.277  LAYER M3  ;
        ANTENNAPARTIALMETALSIDEAREA 96.916  LAYER M2  ;
        ANTENNAPARTIALMETALSIDEAREA 67.374  LAYER M1  ;
        ANTENNADIFFAREA 20.600  LAYER M3  ;
        ANTENNAPARTIALCUTAREA 0.135  LAYER V3  ;
        ANTENNAPARTIALCUTAREA 0.203  LAYER V2  ;
        PORT
        LAYER M3 ;
        RECT  28.870 249.580 29.600 250.000 ;
        LAYER M2 ;
        RECT  28.870 249.580 29.600 250.000 ;
        END
    END CIN
    PIN I
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 80.804  LAYER M2  ;
        ANTENNAPARTIALMETALSIDEAREA 67.374  LAYER M1  ;
        ANTENNAPARTIALMETALSIDEAREA 41.096  LAYER M3  ;
        ANTENNADIFFAREA 0.250  LAYER M3  ;
        ANTENNAPARTIALCUTAREA 0.203  LAYER V2  ;
        ANTENNAPARTIALCUTAREA 0.135  LAYER V3  ;
        ANTENNAGATEAREA 8.100  LAYER M2  ;
        ANTENNAGATEAREA 9.900  LAYER M3  ;
        PORT
        LAYER M3 ;
        RECT  27.840 249.580 28.570 250.000 ;
        LAYER M2 ;
        RECT  27.840 249.580 28.570 250.000 ;
        END
    END I
    PIN VDDO
        DIRECTION INOUT ;
        USE power ;
        PORT
        LAYER M3 ;
        RECT  64.200 192.330 65.000 200.640 ;
        RECT  0.000 201.660 65.000 221.520 ;
        RECT  0.000 222.720 65.000 246.820 ;
        RECT  0.000 192.330 0.800 200.640 ;
        LAYER M2 ;
        RECT  0.000 186.470 65.000 195.650 ;
        LAYER TOP_M ;
        RECT  0.000 195.170 65.000 200.640 ;
        RECT  0.000 201.660 65.000 221.520 ;
        RECT  0.000 222.720 65.000 246.820 ;
        END
    END VDDO
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        PORT
        LAYER M3 ;
        RECT  64.200 163.510 65.000 190.890 ;
        RECT  0.000 163.510 0.800 190.890 ;
        LAYER M2 ;
        RECT  0.000 172.080 65.000 183.060 ;
        LAYER TOP_M ;
        RECT  0.000 163.500 65.000 194.560 ;
        END
    END VDD
    PIN VSSO
        DIRECTION INOUT ;
        USE ground ;
        PORT
        LAYER M3 ;
        RECT  0.000 92.060 65.000 123.250 ;
        RECT  64.200 149.940 65.000 162.610 ;
        RECT  0.000 149.940 0.800 162.610 ;
        LAYER M2 ;
        RECT  0.000 147.040 65.000 154.520 ;
        LAYER TOP_M ;
        RECT  0.000 92.060 65.000 123.250 ;
        RECT  0.000 155.410 65.000 162.610 ;
        END
    END VSSO
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        PORT
        LAYER M3 ;
        RECT  64.200 130.690 65.000 148.880 ;
        RECT  0.000 130.690 0.800 148.880 ;
        LAYER M2 ;
        RECT  0.000 136.310 65.000 146.340 ;
        LAYER TOP_M ;
        RECT  0.000 123.850 65.000 154.560 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  2.000 0.000 63.000 250.000 ;
        RECT  0.000 88.990 65.000 130.360 ;
        RECT  0.000 136.510 65.000 157.550 ;
        RECT  0.315 158.150 64.700 158.460 ;
        RECT  0.300 158.930 64.700 159.230 ;
        RECT  0.300 159.530 64.700 159.830 ;
        RECT  0.300 160.130 64.700 160.430 ;
        RECT  0.300 160.730 64.700 161.030 ;
        RECT  0.300 161.330 64.700 161.630 ;
        RECT  0.300 161.910 64.700 162.190 ;
        RECT  0.300 162.490 64.700 162.770 ;
        RECT  0.300 163.070 64.700 163.350 ;
        RECT  0.300 163.650 64.700 163.950 ;
        RECT  0.300 164.250 64.700 164.550 ;
        RECT  0.300 164.850 64.700 165.150 ;
        RECT  0.300 165.450 64.700 165.750 ;
        RECT  0.300 166.050 64.700 166.350 ;
        RECT  0.300 166.650 64.700 166.960 ;
        RECT  0.300 167.260 64.700 167.560 ;
        RECT  0.300 167.860 64.700 168.160 ;
        RECT  0.000 169.150 65.000 197.240 ;
        RECT  0.600 0.600 64.400 250.000 ;
        RECT  0.000 198.470 65.000 250.000 ;
        LAYER M2 ;
        RECT  1.840 196.420 2.120 249.400 ;
        RECT  63.180 196.430 63.670 249.400 ;
        RECT  0.600 196.440 64.400 245.485 ;
        RECT  26.530 196.440 64.400 248.790 ;
        RECT  0.600 196.440 22.950 249.400 ;
        RECT  26.530 196.440 27.050 249.400 ;
        RECT  31.420 196.440 64.400 249.400 ;
        RECT  14.290 183.720 52.380 185.680 ;
        RECT  0.600 183.850 64.400 185.680 ;
        RECT  54.910 183.850 57.160 185.865 ;
        RECT  46.230 183.720 51.730 185.870 ;
        RECT  18.450 155.160 18.800 171.290 ;
        RECT  19.100 155.140 19.420 171.290 ;
        RECT  49.250 155.125 51.490 171.290 ;
        RECT  52.430 155.295 52.740 171.290 ;
        RECT  53.655 155.035 53.935 171.290 ;
        RECT  56.365 155.280 56.645 171.315 ;
        RECT  57.120 155.300 57.400 171.315 ;
        RECT  57.835 155.130 58.115 171.315 ;
        RECT  0.600 155.310 64.400 171.290 ;
        RECT  56.240 155.310 61.880 171.315 ;
        RECT  53.895 155.310 55.870 171.370 ;
        RECT  3.210 155.310 3.490 171.380 ;
        RECT  34.655 155.310 38.715 171.480 ;
        RECT  39.605 155.310 42.020 171.480 ;
        RECT  2.000 0.000 63.000 60.210 ;
        RECT  0.600 0.600 64.400 60.210 ;
        RECT  0.600 0.600 1.210 135.520 ;
        RECT  0.600 91.020 64.400 135.520 ;
        RECT  4.080 91.020 60.940 135.690 ;
        RECT  62.580 91.020 62.995 135.710 ;
        LAYER M3 ;
        RECT  0.600 247.660 23.220 248.740 ;
        RECT  0.600 247.660 22.900 249.400 ;
        RECT  26.260 247.660 64.400 248.740 ;
        RECT  26.580 247.660 27.000 249.400 ;
        RECT  31.470 247.660 64.400 249.400 ;
        RECT  0.600 124.090 64.400 129.850 ;
        RECT  3.990 123.970 60.900 135.790 ;
        RECT  1.640 124.090 63.600 135.790 ;
        RECT  1.810 124.090 2.830 154.520 ;
        RECT  5.155 123.970 60.900 171.560 ;
        RECT  1.640 155.040 63.600 171.560 ;
        RECT  1.640 183.580 63.600 185.950 ;
        RECT  5.490 124.090 63.600 200.820 ;
        RECT  1.640 196.170 63.600 200.820 ;
        RECT  56.300 123.970 56.580 201.060 ;
        RECT  0.600 0.600 64.400 60.480 ;
        RECT  2.000 0.000 63.000 88.700 ;
        RECT  0.600 0.600 1.480 91.220 ;
        RECT  0.600 90.750 64.400 91.220 ;
        LAYER TOP_M ;
        RECT  0.600 247.690 64.400 248.850 ;
        RECT  0.600 247.690 23.010 249.400 ;
        RECT  26.470 247.690 27.110 249.400 ;
        RECT  31.360 247.690 64.400 249.400 ;
        RECT  2.000 0.000 63.000 91.190 ;
        RECT  0.600 0.600 64.400 91.190 ;
    END
END pt3b01d

MACRO pt3b01
    CLASS PAD ;
    FOREIGN pt3b01 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 65.000 BY 250.000 ;
    SYMMETRY X Y R90 ;
    SITE IOSite_c ;
    PIN PAD
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 55.440  LAYER TOP_M  ;
        ANTENNAPARTIALMETALSIDEAREA 287.938  LAYER M3  ;
        ANTENNAPARTIALMETALSIDEAREA 480.740  LAYER M2  ;
        ANTENNADIFFAREA 2657.280  LAYER TOP_M  ;
        ANTENNADIFFAREA 2657.280  LAYER M3  ;
        ANTENNADIFFAREA 1209.600  LAYER M2  ;
        ANTENNAPARTIALCUTAREA 632.318  LAYER TOP_V  ;
        ANTENNAPARTIALCUTAREA 349.898  LAYER V3  ;
        ANTENNAPARTIALCUTAREA 255.798  LAYER V2  ;
        PORT
        LAYER M3 ;
        RECT  23.740 249.580 25.740 250.000 ;
        LAYER M2 ;
        RECT  2.000 61.000 63.000 90.230 ;
        RECT  23.740 246.275 25.740 250.000 ;
        END
    END PAD
    PIN OEN
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 67.374  LAYER M1  ;
        ANTENNAPARTIALMETALSIDEAREA 80.634  LAYER M2  ;
        ANTENNAPARTIALMETALSIDEAREA 41.679  LAYER M3  ;
        ANTENNADIFFAREA 0.250  LAYER M3  ;
        ANTENNAPARTIALCUTAREA 0.203  LAYER V2  ;
        ANTENNAPARTIALCUTAREA 0.135  LAYER V3  ;
        ANTENNAGATEAREA 8.100  LAYER M2  ;
        ANTENNAGATEAREA 9.900  LAYER M3  ;
        PORT
        LAYER M3 ;
        RECT  29.900 249.580 30.630 250.000 ;
        LAYER M2 ;
        RECT  29.900 249.580 30.630 250.000 ;
        END
    END OEN
    PIN CIN
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 32.277  LAYER M3  ;
        ANTENNAPARTIALMETALSIDEAREA 96.916  LAYER M2  ;
        ANTENNAPARTIALMETALSIDEAREA 67.374  LAYER M1  ;
        ANTENNADIFFAREA 20.600  LAYER M3  ;
        ANTENNAPARTIALCUTAREA 0.135  LAYER V3  ;
        ANTENNAPARTIALCUTAREA 0.203  LAYER V2  ;
        PORT
        LAYER M3 ;
        RECT  28.870 249.580 29.600 250.000 ;
        LAYER M2 ;
        RECT  28.870 249.580 29.600 250.000 ;
        END
    END CIN
    PIN I
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 80.804  LAYER M2  ;
        ANTENNAPARTIALMETALSIDEAREA 67.374  LAYER M1  ;
        ANTENNAPARTIALMETALSIDEAREA 41.096  LAYER M3  ;
        ANTENNADIFFAREA 0.250  LAYER M3  ;
        ANTENNAPARTIALCUTAREA 0.203  LAYER V2  ;
        ANTENNAPARTIALCUTAREA 0.135  LAYER V3  ;
        ANTENNAGATEAREA 8.100  LAYER M2  ;
        ANTENNAGATEAREA 9.900  LAYER M3  ;
        PORT
        LAYER M3 ;
        RECT  27.840 249.580 28.570 250.000 ;
        LAYER M2 ;
        RECT  27.840 249.580 28.570 250.000 ;
        END
    END I
    PIN VDDO
        DIRECTION INOUT ;
        USE power ;
        PORT
        LAYER M3 ;
        RECT  64.200 192.330 65.000 200.640 ;
        RECT  0.000 201.660 65.000 221.520 ;
        RECT  0.000 222.720 65.000 246.820 ;
        RECT  0.000 192.330 0.800 200.640 ;
        LAYER M2 ;
        RECT  0.000 186.470 65.000 195.650 ;
        LAYER TOP_M ;
        RECT  0.000 195.170 65.000 200.640 ;
        RECT  0.000 201.660 65.000 221.520 ;
        RECT  0.000 222.720 65.000 246.820 ;
        END
    END VDDO
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        PORT
        LAYER M3 ;
        RECT  64.200 163.510 65.000 190.890 ;
        RECT  0.000 163.510 0.800 190.890 ;
        LAYER M2 ;
        RECT  0.000 172.080 65.000 183.060 ;
        LAYER TOP_M ;
        RECT  0.000 163.500 65.000 194.560 ;
        END
    END VDD
    PIN VSSO
        DIRECTION INOUT ;
        USE ground ;
        PORT
        LAYER M3 ;
        RECT  0.000 92.060 65.000 123.250 ;
        RECT  64.200 149.940 65.000 162.610 ;
        RECT  0.000 149.940 0.800 162.610 ;
        LAYER M2 ;
        RECT  0.000 147.040 65.000 154.520 ;
        LAYER TOP_M ;
        RECT  0.000 92.060 65.000 123.250 ;
        RECT  0.000 155.410 65.000 162.610 ;
        END
    END VSSO
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        PORT
        LAYER M3 ;
        RECT  64.200 130.690 65.000 148.880 ;
        RECT  0.000 130.690 0.800 148.880 ;
        LAYER M2 ;
        RECT  0.000 136.310 65.000 146.340 ;
        LAYER TOP_M ;
        RECT  0.000 123.850 65.000 154.560 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  2.000 0.000 63.000 250.000 ;
        RECT  0.000 88.990 65.000 130.360 ;
        RECT  0.000 136.510 65.000 157.550 ;
        RECT  0.315 158.150 64.700 158.460 ;
        RECT  0.300 158.930 64.700 159.230 ;
        RECT  0.300 159.530 64.700 159.830 ;
        RECT  0.300 160.130 64.700 160.430 ;
        RECT  0.300 160.730 64.700 161.030 ;
        RECT  0.300 161.330 64.700 161.630 ;
        RECT  0.300 161.910 64.700 162.190 ;
        RECT  0.300 162.490 64.700 162.770 ;
        RECT  0.300 163.070 64.700 163.350 ;
        RECT  0.300 163.650 64.700 163.950 ;
        RECT  0.300 164.250 64.700 164.550 ;
        RECT  0.300 164.850 64.700 165.150 ;
        RECT  0.300 165.450 64.700 165.750 ;
        RECT  0.300 166.050 64.700 166.350 ;
        RECT  0.300 166.650 64.700 166.960 ;
        RECT  0.300 167.260 64.700 167.560 ;
        RECT  0.300 167.860 64.700 168.160 ;
        RECT  0.000 169.150 65.000 197.240 ;
        RECT  0.600 0.600 64.400 250.000 ;
        RECT  0.000 198.470 65.000 250.000 ;
        LAYER M2 ;
        RECT  1.840 196.420 2.120 249.400 ;
        RECT  63.180 196.430 63.670 249.400 ;
        RECT  0.600 196.440 64.400 245.485 ;
        RECT  26.530 196.440 64.400 248.790 ;
        RECT  0.600 196.440 22.950 249.400 ;
        RECT  26.530 196.440 27.050 249.400 ;
        RECT  31.420 196.440 64.400 249.400 ;
        RECT  14.290 183.720 52.380 185.680 ;
        RECT  0.600 183.850 64.400 185.680 ;
        RECT  54.910 183.850 57.160 185.865 ;
        RECT  46.230 183.720 51.730 185.870 ;
        RECT  18.450 155.160 18.800 171.290 ;
        RECT  19.100 155.140 19.420 171.290 ;
        RECT  53.655 155.035 53.935 171.290 ;
        RECT  56.365 155.280 56.645 171.315 ;
        RECT  57.120 155.300 57.400 171.315 ;
        RECT  57.835 155.130 58.115 171.315 ;
        RECT  0.600 155.310 64.400 171.290 ;
        RECT  56.240 155.310 61.880 171.315 ;
        RECT  53.895 155.310 55.870 171.370 ;
        RECT  3.210 155.310 3.490 171.380 ;
        RECT  34.655 155.310 38.715 171.480 ;
        RECT  39.605 155.310 42.020 171.480 ;
        RECT  2.000 0.000 63.000 60.210 ;
        RECT  0.600 0.600 64.400 60.210 ;
        RECT  0.600 0.600 1.210 135.520 ;
        RECT  0.600 91.020 64.400 135.520 ;
        RECT  4.080 91.020 60.940 135.690 ;
        RECT  62.580 91.020 62.995 135.710 ;
        LAYER M3 ;
        RECT  0.600 247.660 23.220 248.740 ;
        RECT  0.600 247.660 22.900 249.400 ;
        RECT  26.260 247.660 64.400 248.740 ;
        RECT  26.580 247.660 27.000 249.400 ;
        RECT  31.470 247.660 64.400 249.400 ;
        RECT  0.600 124.090 64.400 129.850 ;
        RECT  3.990 123.970 60.900 135.790 ;
        RECT  1.640 124.090 63.600 135.790 ;
        RECT  1.810 124.090 2.830 154.520 ;
        RECT  5.155 123.970 60.900 171.560 ;
        RECT  1.640 155.040 63.600 171.560 ;
        RECT  1.640 183.580 63.600 185.950 ;
        RECT  5.490 124.090 63.600 200.820 ;
        RECT  1.640 196.170 63.600 200.820 ;
        RECT  56.300 123.970 56.580 201.060 ;
        RECT  0.600 0.600 64.400 60.480 ;
        RECT  2.000 0.000 63.000 88.700 ;
        RECT  0.600 0.600 1.480 91.220 ;
        RECT  0.600 90.750 64.400 91.220 ;
        LAYER TOP_M ;
        RECT  0.600 247.690 64.400 248.850 ;
        RECT  0.600 247.690 23.010 249.400 ;
        RECT  26.470 247.690 27.110 249.400 ;
        RECT  31.360 247.690 64.400 249.400 ;
        RECT  2.000 0.000 63.000 91.190 ;
        RECT  0.600 0.600 64.400 91.190 ;
    END
END pt3b01

MACRO pc3x13
    CLASS PAD ;
    FOREIGN pc3x13 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 130.000 BY 250.000 ;
    SYMMETRY X Y R90 ;
    SITE IOSite_c ;
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 67.946  LAYER M1  ;
        ANTENNAPARTIALMETALSIDEAREA 36.305  LAYER M3  ;
        ANTENNAPARTIALMETALSIDEAREA 80.846  LAYER M2  ;
        ANTENNADIFFAREA 35.840  LAYER M3  ;
        ANTENNAPARTIALCUTAREA 0.135  LAYER V3  ;
        ANTENNAPARTIALCUTAREA 0.203  LAYER V2  ;
        PORT
        LAYER M3 ;
        RECT  28.870 249.620 29.600 250.000 ;
        LAYER M2 ;
        RECT  28.870 249.620 29.600 250.000 ;
        END
    END Z
    PIN EN
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 80.115  LAYER M2  ;
        ANTENNAPARTIALMETALSIDEAREA 67.946  LAYER M1  ;
        ANTENNAPARTIALMETALSIDEAREA 42.861  LAYER M3  ;
        ANTENNADIFFAREA 2.250  LAYER M3  ;
        ANTENNAPARTIALCUTAREA 0.068  LAYER V2  ;
        ANTENNAPARTIALCUTAREA 0.135  LAYER V3  ;
        ANTENNAGATEAREA 12.060  LAYER M3  ;
        PORT
        LAYER M3 ;
        RECT  29.900 249.620 30.630 250.000 ;
        LAYER M2 ;
        RECT  29.900 249.620 30.630 250.000 ;
        END
    END EN
    PIN XIN
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 55.440  LAYER TOP_M  ;
        ANTENNAPARTIALMETALSIDEAREA 205.937  LAYER M3  ;
        ANTENNAPARTIALMETALSIDEAREA 480.740  LAYER M2  ;
        ANTENNADIFFAREA 2657.280  LAYER TOP_M  ;
        ANTENNADIFFAREA 2657.280  LAYER M3  ;
        ANTENNADIFFAREA 1209.600  LAYER M2  ;
        ANTENNAPARTIALCUTAREA 632.318  LAYER TOP_V  ;
        ANTENNAPARTIALCUTAREA 349.898  LAYER V3  ;
        ANTENNAPARTIALCUTAREA 255.798  LAYER V2  ;
        PORT
        LAYER M2 ;
        RECT  67.000 61.000 128.000 90.230 ;
        END
    END XIN
    PIN XOUT
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 55.440  LAYER TOP_M  ;
        ANTENNAPARTIALMETALSIDEAREA 209.753  LAYER M3  ;
        ANTENNAPARTIALMETALSIDEAREA 480.740  LAYER M2  ;
        ANTENNADIFFAREA 2524.080  LAYER TOP_M  ;
        ANTENNADIFFAREA 2524.080  LAYER M3  ;
        ANTENNADIFFAREA 1076.400  LAYER M2  ;
        ANTENNAPARTIALCUTAREA 632.318  LAYER TOP_V  ;
        ANTENNAPARTIALCUTAREA 352.264  LAYER V3  ;
        ANTENNAPARTIALCUTAREA 255.798  LAYER V2  ;
        PORT
        LAYER M2 ;
        RECT  2.000 61.000 63.000 90.230 ;
        END
    END XOUT
    PIN VDDO
        DIRECTION INOUT ;
        USE power ;
        PORT
        LAYER TOP_M ;
        RECT  0.000 195.170 130.000 200.640 ;
        RECT  0.000 201.660 130.000 221.520 ;
        RECT  0.000 222.720 130.000 246.820 ;
        LAYER M3 ;
        RECT  129.200 192.330 130.000 200.640 ;
        RECT  0.000 222.720 130.000 246.820 ;
        RECT  0.000 201.660 130.000 221.520 ;
        RECT  0.000 192.330 0.800 200.640 ;
        LAYER M2 ;
        RECT  62.630 186.470 130.000 195.650 ;
        RECT  0.000 186.470 130.000 190.060 ;
        RECT  0.000 186.470 2.745 195.650 ;
        END
    END VDDO
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        PORT
        LAYER TOP_M ;
        RECT  0.000 163.500 130.000 194.560 ;
        LAYER M3 ;
        RECT  129.200 163.510 130.000 190.890 ;
        RECT  0.000 163.510 0.800 190.890 ;
        LAYER M2 ;
        RECT  124.230 172.080 130.000 183.060 ;
        RECT  0.000 175.005 130.000 179.440 ;
        RECT  96.040 172.080 130.000 179.440 ;
        RECT  0.000 175.005 94.540 183.060 ;
        RECT  0.000 172.080 72.710 183.060 ;
        END
    END VDD
    PIN VSSO
        DIRECTION INOUT ;
        USE ground ;
        PORT
        LAYER TOP_M ;
        RECT  0.000 92.060 130.000 123.250 ;
        RECT  0.000 155.410 130.000 162.610 ;
        LAYER M3 ;
        RECT  63.650 92.060 130.000 123.250 ;
        RECT  0.000 92.060 130.000 122.010 ;
        RECT  0.000 92.060 2.975 123.250 ;
        RECT  129.200 149.940 130.000 162.610 ;
        RECT  0.000 149.940 0.800 162.610 ;
        LAYER M2 ;
        RECT  0.000 147.040 130.000 154.520 ;
        END
    END VSSO
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        PORT
        LAYER TOP_M ;
        RECT  0.000 123.850 130.000 154.560 ;
        LAYER M3 ;
        RECT  129.200 130.690 130.000 148.880 ;
        RECT  0.000 130.690 0.800 148.880 ;
        LAYER M2 ;
        RECT  0.000 136.310 130.000 146.340 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  2.000 0.000 63.000 250.000 ;
        RECT  67.000 0.000 128.000 250.000 ;
        RECT  0.000 88.990 130.000 130.360 ;
        RECT  0.000 136.510 130.000 157.550 ;
        RECT  0.300 158.930 129.700 159.230 ;
        RECT  0.300 159.530 129.700 159.830 ;
        RECT  0.300 160.130 129.700 160.430 ;
        RECT  0.300 160.730 129.700 161.030 ;
        RECT  0.300 161.330 129.700 161.630 ;
        RECT  0.300 161.910 129.700 162.190 ;
        RECT  0.300 162.490 129.700 162.770 ;
        RECT  0.300 163.070 129.700 163.350 ;
        RECT  0.300 163.650 129.700 163.950 ;
        RECT  0.300 164.250 129.700 164.550 ;
        RECT  0.300 164.850 129.700 165.150 ;
        RECT  0.300 165.450 129.700 165.750 ;
        RECT  0.300 166.050 129.700 166.350 ;
        RECT  0.300 166.650 129.700 166.960 ;
        RECT  0.300 167.260 129.700 167.560 ;
        RECT  0.300 167.860 129.700 168.160 ;
        RECT  0.600 0.600 129.400 250.000 ;
        RECT  0.000 198.470 130.000 250.000 ;
        LAYER M2 ;
        RECT  6.800 190.840 8.920 249.400 ;
        RECT  3.535 190.850 61.840 248.830 ;
        RECT  0.600 196.440 28.080 249.400 ;
        RECT  31.420 196.440 129.400 249.400 ;
        RECT  89.710 183.845 94.390 185.680 ;
        RECT  95.330 180.230 123.440 185.680 ;
        RECT  0.600 183.850 129.400 185.680 ;
        RECT  12.220 183.850 14.320 185.700 ;
        RECT  118.395 183.660 123.505 185.865 ;
        RECT  2.905 155.015 14.445 171.290 ;
        RECT  27.410 155.260 27.880 171.290 ;
        RECT  33.690 155.120 34.010 171.430 ;
        RECT  52.335 155.175 52.905 171.290 ;
        RECT  56.955 155.160 57.370 171.290 ;
        RECT  57.975 155.000 58.330 171.290 ;
        RECT  60.405 155.290 60.905 171.290 ;
        RECT  69.685 155.235 69.995 171.290 ;
        RECT  70.730 155.200 71.040 171.290 ;
        RECT  0.600 155.310 129.400 171.290 ;
        RECT  127.450 154.990 128.380 171.380 ;
        RECT  73.500 155.310 128.380 171.380 ;
        RECT  30.410 155.310 34.090 171.430 ;
        RECT  34.410 155.310 34.730 171.480 ;
        RECT  73.500 155.310 95.250 174.215 ;
        RECT  74.570 155.310 94.960 174.455 ;
        RECT  2.000 0.000 63.000 60.210 ;
        RECT  67.000 0.000 128.000 60.210 ;
        RECT  0.600 0.600 129.400 60.210 ;
        RECT  63.790 0.600 66.210 135.520 ;
        RECT  0.600 91.020 129.400 135.520 ;
        RECT  4.070 91.020 60.930 135.690 ;
        RECT  69.000 91.020 125.860 135.690 ;
        RECT  2.905 91.020 3.470 135.710 ;
        LAYER M3 ;
        RECT  0.600 247.660 129.400 248.780 ;
        RECT  0.600 247.660 28.030 249.400 ;
        RECT  31.470 247.660 129.400 249.400 ;
        RECT  3.815 122.850 62.810 200.820 ;
        RECT  68.960 124.070 126.190 171.560 ;
        RECT  0.600 124.090 129.400 129.850 ;
        RECT  1.400 124.090 128.360 135.790 ;
        RECT  127.170 124.090 128.190 154.520 ;
        RECT  1.400 124.090 126.190 160.480 ;
        RECT  1.640 155.040 128.360 171.560 ;
        RECT  1.640 183.580 128.360 185.950 ;
        RECT  2.745 124.090 124.660 200.820 ;
        RECT  1.640 196.170 128.360 200.820 ;
        RECT  2.745 124.090 3.115 200.840 ;
        RECT  66.190 124.090 117.430 221.880 ;
        RECT  0.600 0.600 129.400 60.480 ;
        RECT  2.000 0.000 63.000 88.700 ;
        RECT  67.000 0.000 128.000 88.700 ;
        RECT  63.520 0.600 66.480 91.220 ;
        RECT  0.600 90.750 129.400 91.220 ;
        LAYER TOP_M ;
        RECT  0.600 247.690 129.400 248.890 ;
        RECT  0.600 247.690 28.140 249.400 ;
        RECT  31.360 247.690 129.400 249.400 ;
        RECT  2.000 0.000 63.000 91.190 ;
        RECT  67.000 0.000 128.000 91.190 ;
        RECT  0.600 0.600 129.400 91.190 ;
    END
END pc3x13

MACRO pc3x12
    CLASS PAD ;
    FOREIGN pc3x12 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 130.000 BY 250.000 ;
    SYMMETRY X Y R90 ;
    SITE IOSite_c ;
    PIN XIN
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 55.440  LAYER TOP_M  ;
        ANTENNAPARTIALMETALSIDEAREA 205.937  LAYER M3  ;
        ANTENNAPARTIALMETALSIDEAREA 480.740  LAYER M2  ;
        ANTENNADIFFAREA 2657.280  LAYER TOP_M  ;
        ANTENNADIFFAREA 2657.280  LAYER M3  ;
        ANTENNADIFFAREA 1209.600  LAYER M2  ;
        ANTENNAPARTIALCUTAREA 632.318  LAYER TOP_V  ;
        ANTENNAPARTIALCUTAREA 349.898  LAYER V3  ;
        ANTENNAPARTIALCUTAREA 255.798  LAYER V2  ;
        PORT
        LAYER M2 ;
        RECT  67.000 61.000 128.000 90.230 ;
        END
    END XIN
    PIN XOUT
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 55.440  LAYER TOP_M  ;
        ANTENNAPARTIALMETALSIDEAREA 209.753  LAYER M3  ;
        ANTENNAPARTIALMETALSIDEAREA 480.740  LAYER M2  ;
        ANTENNADIFFAREA 2580.480  LAYER TOP_M  ;
        ANTENNADIFFAREA 2580.480  LAYER M3  ;
        ANTENNADIFFAREA 1132.800  LAYER M2  ;
        ANTENNAPARTIALCUTAREA 632.318  LAYER TOP_V  ;
        ANTENNAPARTIALCUTAREA 352.264  LAYER V3  ;
        ANTENNAPARTIALCUTAREA 255.798  LAYER V2  ;
        PORT
        LAYER M2 ;
        RECT  2.000 61.000 63.000 90.230 ;
        END
    END XOUT
    PIN EN
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 67.946  LAYER M1  ;
        ANTENNAPARTIALMETALSIDEAREA 42.861  LAYER M3  ;
        ANTENNAPARTIALMETALSIDEAREA 80.115  LAYER M2  ;
        ANTENNADIFFAREA 2.250  LAYER M3  ;
        ANTENNAPARTIALCUTAREA 0.135  LAYER V3  ;
        ANTENNAPARTIALCUTAREA 0.068  LAYER V2  ;
        ANTENNAGATEAREA 12.060  LAYER M3  ;
        PORT
        LAYER M3 ;
        RECT  29.900 249.620 30.630 250.000 ;
        LAYER M2 ;
        RECT  29.900 249.620 30.630 250.000 ;
        END
    END EN
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 67.946  LAYER M1  ;
        ANTENNAPARTIALMETALSIDEAREA 36.305  LAYER M3  ;
        ANTENNAPARTIALMETALSIDEAREA 80.846  LAYER M2  ;
        ANTENNADIFFAREA 35.840  LAYER M3  ;
        ANTENNAPARTIALCUTAREA 0.135  LAYER V3  ;
        ANTENNAPARTIALCUTAREA 0.203  LAYER V2  ;
        PORT
        LAYER M3 ;
        RECT  28.870 249.620 29.600 250.000 ;
        LAYER M2 ;
        RECT  28.870 249.620 29.600 250.000 ;
        END
    END Z
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        PORT
        LAYER M3 ;
        RECT  129.200 130.690 130.000 148.880 ;
        RECT  0.000 130.690 0.800 148.880 ;
        LAYER TOP_M ;
        RECT  0.000 123.850 130.000 154.560 ;
        LAYER M2 ;
        RECT  0.000 136.310 130.000 146.340 ;
        END
    END VSS
    PIN VSSO
        DIRECTION INOUT ;
        USE ground ;
        PORT
        LAYER M3 ;
        RECT  63.650 92.060 130.000 123.250 ;
        RECT  0.000 92.060 130.000 122.430 ;
        RECT  0.000 92.060 2.975 123.250 ;
        RECT  129.200 149.940 130.000 162.610 ;
        RECT  0.000 149.940 0.800 162.610 ;
        LAYER TOP_M ;
        RECT  0.000 92.060 130.000 123.250 ;
        RECT  0.000 155.410 130.000 162.610 ;
        LAYER M2 ;
        RECT  0.000 147.040 130.000 154.520 ;
        END
    END VSSO
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        PORT
        LAYER M3 ;
        RECT  129.200 163.510 130.000 190.890 ;
        RECT  0.000 163.510 0.800 190.890 ;
        LAYER TOP_M ;
        RECT  0.000 163.500 130.000 194.560 ;
        LAYER M2 ;
        RECT  124.230 172.080 130.000 183.060 ;
        RECT  0.000 175.005 130.000 179.440 ;
        RECT  96.040 172.080 130.000 179.440 ;
        RECT  0.000 175.005 94.540 183.060 ;
        RECT  0.000 172.080 72.710 183.060 ;
        END
    END VDD
    PIN VDDO
        DIRECTION INOUT ;
        USE power ;
        PORT
        LAYER M3 ;
        RECT  129.200 192.330 130.000 200.640 ;
        RECT  0.000 222.720 130.000 246.820 ;
        RECT  0.000 201.660 130.000 221.520 ;
        RECT  0.000 192.330 0.800 200.640 ;
        LAYER TOP_M ;
        RECT  0.000 195.170 130.000 200.640 ;
        RECT  0.000 201.660 130.000 221.520 ;
        RECT  0.000 222.720 130.000 246.820 ;
        LAYER M2 ;
        RECT  62.630 186.470 130.000 195.650 ;
        RECT  0.000 186.470 130.000 190.060 ;
        RECT  0.000 186.470 2.745 195.650 ;
        END
    END VDDO
    OBS
        LAYER M1 ;
        RECT  2.000 0.000 63.000 250.000 ;
        RECT  67.000 0.000 128.000 250.000 ;
        RECT  0.000 88.990 130.000 130.360 ;
        RECT  0.000 136.510 130.000 157.550 ;
        RECT  0.300 158.930 129.700 159.230 ;
        RECT  0.300 159.530 129.700 159.830 ;
        RECT  0.300 160.130 129.700 160.430 ;
        RECT  0.300 160.730 129.700 161.030 ;
        RECT  0.300 161.330 129.700 161.630 ;
        RECT  0.300 161.910 129.700 162.190 ;
        RECT  0.300 162.490 129.700 162.770 ;
        RECT  0.300 163.070 129.700 163.350 ;
        RECT  0.300 163.650 129.700 163.950 ;
        RECT  0.300 164.250 129.700 164.550 ;
        RECT  0.300 164.850 129.700 165.150 ;
        RECT  0.300 165.450 129.700 165.750 ;
        RECT  0.300 166.050 129.700 166.350 ;
        RECT  0.300 166.650 129.700 166.960 ;
        RECT  0.300 167.260 129.700 167.560 ;
        RECT  0.300 167.860 129.700 168.160 ;
        RECT  0.600 0.600 129.400 250.000 ;
        RECT  0.000 198.470 130.000 250.000 ;
        LAYER M2 ;
        RECT  6.800 190.840 8.920 249.400 ;
        RECT  3.535 190.850 61.840 248.830 ;
        RECT  0.600 196.440 28.080 249.400 ;
        RECT  31.420 196.440 129.400 249.400 ;
        RECT  89.710 183.845 94.390 185.680 ;
        RECT  95.330 180.230 123.440 185.680 ;
        RECT  0.600 183.850 129.400 185.680 ;
        RECT  12.220 183.850 14.320 185.700 ;
        RECT  118.395 183.660 123.505 185.865 ;
        RECT  2.905 155.015 14.445 171.290 ;
        RECT  27.415 155.260 27.885 171.290 ;
        RECT  33.695 155.120 34.015 171.430 ;
        RECT  52.355 155.175 52.925 171.290 ;
        RECT  56.975 155.160 57.390 171.290 ;
        RECT  57.995 155.000 58.350 171.290 ;
        RECT  60.425 155.290 60.925 171.290 ;
        RECT  69.685 155.235 69.995 171.290 ;
        RECT  70.730 155.200 71.040 171.290 ;
        RECT  0.600 155.310 129.400 171.290 ;
        RECT  127.450 154.990 128.380 171.380 ;
        RECT  73.500 155.310 128.380 171.380 ;
        RECT  30.415 155.310 34.095 171.430 ;
        RECT  34.415 155.310 34.735 171.480 ;
        RECT  73.500 155.310 95.250 174.215 ;
        RECT  74.570 155.310 94.960 174.455 ;
        RECT  2.000 0.000 63.000 60.210 ;
        RECT  67.000 0.000 128.000 60.210 ;
        RECT  0.600 0.600 129.400 60.210 ;
        RECT  63.790 0.600 66.210 135.520 ;
        RECT  0.600 91.020 129.400 135.520 ;
        RECT  4.070 91.020 60.930 135.690 ;
        RECT  69.000 91.020 125.860 135.690 ;
        RECT  2.905 91.020 3.470 135.710 ;
        LAYER M3 ;
        RECT  0.600 247.660 129.400 248.780 ;
        RECT  0.600 247.660 28.030 249.400 ;
        RECT  31.470 247.660 129.400 249.400 ;
        RECT  4.125 123.030 60.870 200.820 ;
        RECT  3.815 123.270 62.810 200.820 ;
        RECT  68.960 124.070 126.190 171.560 ;
        RECT  0.600 124.090 129.400 129.850 ;
        RECT  1.400 124.090 128.360 135.790 ;
        RECT  127.170 124.090 128.190 154.520 ;
        RECT  1.400 124.090 126.190 160.515 ;
        RECT  1.640 155.040 128.360 171.560 ;
        RECT  1.640 183.580 128.360 185.950 ;
        RECT  2.725 124.090 124.660 200.820 ;
        RECT  1.640 196.170 128.360 200.820 ;
        RECT  10.390 123.030 10.790 200.900 ;
        RECT  66.190 124.090 117.430 221.880 ;
        RECT  0.600 0.600 129.400 60.480 ;
        RECT  2.000 0.000 63.000 88.700 ;
        RECT  67.000 0.000 128.000 88.700 ;
        RECT  63.520 0.600 66.480 91.220 ;
        RECT  0.600 90.750 129.400 91.220 ;
        LAYER TOP_M ;
        RECT  0.600 247.690 129.400 248.890 ;
        RECT  0.600 247.690 28.140 249.400 ;
        RECT  31.360 247.690 129.400 249.400 ;
        RECT  2.000 0.000 63.000 91.190 ;
        RECT  67.000 0.000 128.000 91.190 ;
        RECT  0.600 0.600 129.400 91.190 ;
    END
END pc3x12

MACRO pc3x11
    CLASS PAD ;
    FOREIGN pc3x11 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 130.000 BY 250.000 ;
    SYMMETRY X Y R90 ;
    SITE IOSite_c ;
    PIN EN
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 80.115  LAYER M2  ;
        ANTENNAPARTIALMETALSIDEAREA 67.946  LAYER M1  ;
        ANTENNAPARTIALMETALSIDEAREA 42.861  LAYER M3  ;
        ANTENNADIFFAREA 2.250  LAYER M3  ;
        ANTENNAPARTIALCUTAREA 0.135  LAYER V3  ;
        ANTENNAPARTIALCUTAREA 0.068  LAYER V2  ;
        ANTENNAGATEAREA 12.060  LAYER M3  ;
        PORT
        LAYER M3 ;
        RECT  29.900 249.620 30.630 250.000 ;
        LAYER M2 ;
        RECT  29.900 249.620 30.630 250.000 ;
        END
    END EN
    PIN Z
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 80.846  LAYER M2  ;
        ANTENNAPARTIALMETALSIDEAREA 67.946  LAYER M1  ;
        ANTENNAPARTIALMETALSIDEAREA 36.305  LAYER M3  ;
        ANTENNADIFFAREA 35.840  LAYER M3  ;
        ANTENNAPARTIALCUTAREA 0.203  LAYER V2  ;
        ANTENNAPARTIALCUTAREA 0.135  LAYER V3  ;
        PORT
        LAYER M3 ;
        RECT  28.870 249.620 29.600 250.000 ;
        LAYER M2 ;
        RECT  28.870 249.620 29.600 250.000 ;
        END
    END Z
    PIN XOUT
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 55.440  LAYER TOP_M  ;
        ANTENNAPARTIALMETALSIDEAREA 209.753  LAYER M3  ;
        ANTENNAPARTIALMETALSIDEAREA 480.740  LAYER M2  ;
        ANTENNADIFFAREA 2636.880  LAYER TOP_M  ;
        ANTENNADIFFAREA 2636.880  LAYER M3  ;
        ANTENNADIFFAREA 1189.200  LAYER M2  ;
        ANTENNAPARTIALCUTAREA 632.318  LAYER TOP_V  ;
        ANTENNAPARTIALCUTAREA 352.264  LAYER V3  ;
        ANTENNAPARTIALCUTAREA 255.798  LAYER V2  ;
        PORT
        LAYER M2 ;
        RECT  2.000 61.000 63.000 90.230 ;
        END
    END XOUT
    PIN XIN
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 55.440  LAYER TOP_M  ;
        ANTENNAPARTIALMETALSIDEAREA 205.937  LAYER M3  ;
        ANTENNAPARTIALMETALSIDEAREA 480.740  LAYER M2  ;
        ANTENNADIFFAREA 2657.280  LAYER TOP_M  ;
        ANTENNADIFFAREA 2657.280  LAYER M3  ;
        ANTENNADIFFAREA 1209.600  LAYER M2  ;
        ANTENNAPARTIALCUTAREA 632.318  LAYER TOP_V  ;
        ANTENNAPARTIALCUTAREA 349.898  LAYER V3  ;
        ANTENNAPARTIALCUTAREA 255.798  LAYER V2  ;
        PORT
        LAYER M2 ;
        RECT  67.000 61.000 128.000 90.230 ;
        END
    END XIN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        PORT
        LAYER M3 ;
        RECT  129.200 130.690 130.000 148.880 ;
        RECT  0.000 130.690 0.800 148.880 ;
        LAYER TOP_M ;
        RECT  0.000 123.850 130.000 154.560 ;
        LAYER M2 ;
        RECT  0.000 136.310 130.000 146.340 ;
        END
    END VSS
    PIN VSSO
        DIRECTION INOUT ;
        USE ground ;
        PORT
        LAYER M3 ;
        RECT  63.650 92.060 130.000 123.250 ;
        RECT  0.000 92.060 130.000 122.010 ;
        RECT  0.000 92.060 2.975 123.250 ;
        RECT  129.200 149.940 130.000 162.610 ;
        RECT  0.000 149.940 0.800 162.610 ;
        LAYER TOP_M ;
        RECT  0.000 92.060 130.000 123.250 ;
        RECT  0.000 155.410 130.000 162.610 ;
        LAYER M2 ;
        RECT  0.000 147.040 130.000 154.520 ;
        END
    END VSSO
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        PORT
        LAYER M3 ;
        RECT  129.200 163.510 130.000 190.890 ;
        RECT  0.000 163.510 0.800 190.890 ;
        LAYER TOP_M ;
        RECT  0.000 163.500 130.000 194.560 ;
        LAYER M2 ;
        RECT  124.230 172.080 130.000 183.060 ;
        RECT  0.000 175.005 130.000 179.440 ;
        RECT  96.040 172.080 130.000 179.440 ;
        RECT  0.000 175.005 94.540 183.060 ;
        RECT  0.000 172.080 72.710 183.060 ;
        END
    END VDD
    PIN VDDO
        DIRECTION INOUT ;
        USE power ;
        PORT
        LAYER M3 ;
        RECT  129.200 192.330 130.000 200.640 ;
        RECT  0.000 222.720 130.000 246.820 ;
        RECT  0.000 201.660 130.000 221.520 ;
        RECT  0.000 192.330 0.800 200.640 ;
        LAYER TOP_M ;
        RECT  0.000 195.170 130.000 200.640 ;
        RECT  0.000 201.660 130.000 221.520 ;
        RECT  0.000 222.720 130.000 246.820 ;
        LAYER M2 ;
        RECT  62.630 186.470 130.000 195.650 ;
        RECT  0.000 186.470 130.000 190.060 ;
        RECT  0.000 186.470 2.745 195.650 ;
        END
    END VDDO
    OBS
        LAYER M1 ;
        RECT  2.000 0.000 63.000 250.000 ;
        RECT  67.000 0.000 128.000 250.000 ;
        RECT  0.000 88.990 130.000 130.360 ;
        RECT  0.000 136.510 130.000 157.550 ;
        RECT  0.300 158.930 129.700 159.230 ;
        RECT  0.300 159.530 129.700 159.830 ;
        RECT  0.300 160.130 129.700 160.430 ;
        RECT  0.300 160.730 129.700 161.030 ;
        RECT  0.300 161.330 129.700 161.630 ;
        RECT  0.300 161.910 129.700 162.190 ;
        RECT  0.300 162.490 129.700 162.770 ;
        RECT  0.300 163.070 129.700 163.350 ;
        RECT  0.300 163.650 129.700 163.950 ;
        RECT  0.300 164.250 129.700 164.550 ;
        RECT  0.300 164.850 129.700 165.150 ;
        RECT  0.300 165.450 129.700 165.750 ;
        RECT  0.300 166.050 129.700 166.350 ;
        RECT  0.300 166.650 129.700 166.960 ;
        RECT  0.300 167.260 129.700 167.560 ;
        RECT  0.300 167.860 129.700 168.160 ;
        RECT  0.600 0.600 129.400 250.000 ;
        RECT  0.000 198.470 130.000 250.000 ;
        LAYER M2 ;
        RECT  6.800 190.840 8.920 249.400 ;
        RECT  3.535 190.850 61.840 248.830 ;
        RECT  0.600 196.440 28.080 249.400 ;
        RECT  31.420 196.440 129.400 249.400 ;
        RECT  89.710 183.845 94.390 185.680 ;
        RECT  95.330 180.230 123.440 185.680 ;
        RECT  0.600 183.850 129.400 185.680 ;
        RECT  12.220 183.850 14.320 185.700 ;
        RECT  118.395 183.660 123.505 185.865 ;
        RECT  2.905 155.015 14.445 171.290 ;
        RECT  27.415 155.260 27.885 171.290 ;
        RECT  33.695 155.120 34.015 171.430 ;
        RECT  52.335 155.175 52.905 171.290 ;
        RECT  56.955 155.160 57.370 171.290 ;
        RECT  57.975 155.000 58.330 171.290 ;
        RECT  60.405 155.290 60.905 171.290 ;
        RECT  69.685 155.235 69.995 171.290 ;
        RECT  70.730 155.200 71.040 171.290 ;
        RECT  0.600 155.310 129.400 171.290 ;
        RECT  127.450 154.990 128.380 171.380 ;
        RECT  73.500 155.310 128.380 171.380 ;
        RECT  30.415 155.310 34.095 171.430 ;
        RECT  34.415 155.310 34.735 171.480 ;
        RECT  73.500 155.310 95.250 174.215 ;
        RECT  74.570 155.310 94.960 174.455 ;
        RECT  2.000 0.000 63.000 60.210 ;
        RECT  67.000 0.000 128.000 60.210 ;
        RECT  0.600 0.600 129.400 60.210 ;
        RECT  63.790 0.600 66.210 135.520 ;
        RECT  0.600 91.020 129.400 135.520 ;
        RECT  4.070 91.020 60.930 135.690 ;
        RECT  69.000 91.020 125.860 135.690 ;
        RECT  2.905 91.020 3.470 135.710 ;
        LAYER M3 ;
        RECT  0.600 247.660 129.400 248.780 ;
        RECT  0.600 247.660 28.030 249.400 ;
        RECT  31.470 247.660 129.400 249.400 ;
        RECT  3.815 122.850 62.810 200.820 ;
        RECT  68.960 124.070 126.190 171.560 ;
        RECT  0.600 124.090 129.400 129.850 ;
        RECT  1.400 124.090 128.360 135.790 ;
        RECT  127.170 124.090 128.190 154.520 ;
        RECT  1.400 124.090 126.190 160.480 ;
        RECT  1.640 155.040 128.360 171.560 ;
        RECT  1.640 183.580 128.360 185.950 ;
        RECT  2.670 124.090 124.660 200.820 ;
        RECT  1.640 196.170 128.360 200.820 ;
        RECT  66.190 124.090 117.430 221.880 ;
        RECT  0.600 0.600 129.400 60.480 ;
        RECT  2.000 0.000 63.000 88.700 ;
        RECT  67.000 0.000 128.000 88.700 ;
        RECT  63.520 0.600 66.480 91.220 ;
        RECT  0.600 90.750 129.400 91.220 ;
        LAYER TOP_M ;
        RECT  0.600 247.690 129.400 248.890 ;
        RECT  0.600 247.690 28.140 249.400 ;
        RECT  31.360 247.690 129.400 249.400 ;
        RECT  2.000 0.000 63.000 91.190 ;
        RECT  67.000 0.000 128.000 91.190 ;
        RECT  0.600 0.600 129.400 91.190 ;
    END
END pc3x11

MACRO pc3t05u
    CLASS PAD ;
    FOREIGN pc3t05u 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 65.000 BY 250.000 ;
    SYMMETRY X Y R90 ;
    SITE IOSite_c ;
    PIN PAD
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 55.440  LAYER TOP_M  ;
        ANTENNAPARTIALMETALSIDEAREA 287.938  LAYER M3  ;
        ANTENNAPARTIALMETALSIDEAREA 480.740  LAYER M2  ;
        ANTENNADIFFAREA 2657.280  LAYER TOP_M  ;
        ANTENNADIFFAREA 2657.280  LAYER M3  ;
        ANTENNADIFFAREA 1209.600  LAYER M2  ;
        ANTENNAPARTIALCUTAREA 632.318  LAYER TOP_V  ;
        ANTENNAPARTIALCUTAREA 349.898  LAYER V3  ;
        ANTENNAPARTIALCUTAREA 255.798  LAYER V2  ;
        PORT
        LAYER M3 ;
        RECT  23.740 249.580 25.740 250.000 ;
        LAYER M2 ;
        RECT  2.000 61.000 63.000 90.230 ;
        RECT  23.740 246.275 25.740 250.000 ;
        END
    END PAD
    PIN OEN
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 81.726  LAYER M2  ;
        ANTENNAPARTIALMETALSIDEAREA 67.374  LAYER M1  ;
        ANTENNAPARTIALMETALSIDEAREA 41.679  LAYER M3  ;
        ANTENNADIFFAREA 0.250  LAYER M3  ;
        ANTENNAPARTIALCUTAREA 0.135  LAYER V3  ;
        ANTENNAPARTIALCUTAREA 0.203  LAYER V2  ;
        ANTENNAGATEAREA 8.100  LAYER M2  ;
        ANTENNAGATEAREA 9.900  LAYER M3  ;
        PORT
        LAYER M3 ;
        RECT  28.870 249.580 29.600 250.000 ;
        LAYER M2 ;
        RECT  28.870 249.580 29.600 250.000 ;
        END
    END OEN
    PIN I
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 67.374  LAYER M1  ;
        ANTENNAPARTIALMETALSIDEAREA 80.804  LAYER M2  ;
        ANTENNAPARTIALMETALSIDEAREA 41.096  LAYER M3  ;
        ANTENNADIFFAREA 0.250  LAYER M3  ;
        ANTENNAPARTIALCUTAREA 0.270  LAYER V2  ;
        ANTENNAPARTIALCUTAREA 0.135  LAYER V3  ;
        ANTENNAGATEAREA 18.900  LAYER M2  ;
        ANTENNAGATEAREA 20.700  LAYER M3  ;
        PORT
        LAYER M3 ;
        RECT  27.840 249.580 28.570 250.000 ;
        LAYER M2 ;
        RECT  27.840 249.580 28.570 250.000 ;
        END
    END I
    PIN VDDO
        DIRECTION INOUT ;
        USE power ;
        PORT
        LAYER M3 ;
        RECT  64.200 192.330 65.000 200.640 ;
        RECT  0.000 201.660 65.000 221.520 ;
        RECT  0.000 222.720 65.000 246.820 ;
        RECT  0.000 192.330 0.800 200.640 ;
        LAYER M2 ;
        RECT  0.000 186.470 65.000 195.650 ;
        LAYER TOP_M ;
        RECT  0.000 195.170 65.000 200.640 ;
        RECT  0.000 201.660 65.000 221.520 ;
        RECT  0.000 222.720 65.000 246.820 ;
        END
    END VDDO
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        PORT
        LAYER M3 ;
        RECT  64.200 163.510 65.000 190.890 ;
        RECT  0.000 163.510 0.800 190.890 ;
        LAYER M2 ;
        RECT  0.000 172.080 65.000 183.060 ;
        LAYER TOP_M ;
        RECT  0.000 163.500 65.000 194.560 ;
        END
    END VDD
    PIN VSSO
        DIRECTION INOUT ;
        USE ground ;
        PORT
        LAYER M3 ;
        RECT  0.000 92.060 65.000 123.250 ;
        RECT  64.200 149.940 65.000 162.610 ;
        RECT  0.000 149.940 0.800 162.610 ;
        LAYER M2 ;
        RECT  0.000 147.040 65.000 154.520 ;
        LAYER TOP_M ;
        RECT  0.000 92.060 65.000 123.250 ;
        RECT  0.000 155.410 65.000 162.610 ;
        END
    END VSSO
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        PORT
        LAYER M3 ;
        RECT  64.200 130.690 65.000 148.880 ;
        RECT  0.000 130.690 0.800 148.880 ;
        LAYER M2 ;
        RECT  0.000 136.310 65.000 146.340 ;
        LAYER TOP_M ;
        RECT  0.000 123.850 65.000 154.560 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  2.000 0.000 63.000 250.000 ;
        RECT  0.000 88.990 65.000 130.360 ;
        RECT  0.000 136.510 65.000 157.550 ;
        RECT  0.315 158.150 64.700 158.460 ;
        RECT  0.300 158.930 64.700 159.230 ;
        RECT  0.300 159.530 64.700 159.830 ;
        RECT  0.300 160.130 64.700 160.430 ;
        RECT  0.300 160.730 64.700 161.030 ;
        RECT  0.300 161.330 64.700 161.630 ;
        RECT  0.300 161.910 64.700 162.190 ;
        RECT  0.300 162.490 64.700 162.770 ;
        RECT  0.300 163.070 64.700 163.350 ;
        RECT  0.300 163.650 64.700 163.950 ;
        RECT  0.300 164.250 64.700 164.550 ;
        RECT  0.300 164.850 64.700 165.150 ;
        RECT  0.300 165.450 64.700 165.750 ;
        RECT  0.300 166.050 64.700 166.350 ;
        RECT  0.300 166.650 64.700 166.960 ;
        RECT  0.300 167.260 64.700 167.560 ;
        RECT  0.300 167.860 64.700 168.160 ;
        RECT  0.000 169.150 65.000 197.240 ;
        RECT  0.600 0.600 64.400 250.000 ;
        RECT  0.000 198.470 65.000 250.000 ;
        LAYER M2 ;
        RECT  63.180 196.430 63.670 249.400 ;
        RECT  0.600 196.440 64.400 245.485 ;
        RECT  26.530 196.440 64.400 248.790 ;
        RECT  0.600 196.440 22.950 249.400 ;
        RECT  26.530 196.440 27.050 249.400 ;
        RECT  30.390 196.440 64.400 249.400 ;
        RECT  0.600 183.850 64.400 185.680 ;
        RECT  46.230 183.850 51.730 185.870 ;
        RECT  4.480 154.920 7.530 171.290 ;
        RECT  8.170 155.125 8.490 171.290 ;
        RECT  21.210 155.160 21.560 171.290 ;
        RECT  21.860 155.140 22.180 171.290 ;
        RECT  31.895 155.120 35.765 171.290 ;
        RECT  53.655 155.035 53.935 171.290 ;
        RECT  56.365 155.280 56.645 171.290 ;
        RECT  57.120 155.300 57.400 171.290 ;
        RECT  57.835 155.130 58.115 171.290 ;
        RECT  0.600 155.310 64.400 171.290 ;
        RECT  53.895 155.310 55.870 171.370 ;
        RECT  3.170 155.310 3.450 171.380 ;
        RECT  34.655 155.310 38.715 171.480 ;
        RECT  39.605 155.310 42.020 171.480 ;
        RECT  2.000 0.000 63.000 60.210 ;
        RECT  0.600 0.600 64.400 60.210 ;
        RECT  0.600 0.600 1.210 135.520 ;
        RECT  0.600 91.020 64.400 135.520 ;
        RECT  4.080 91.020 60.940 135.690 ;
        RECT  62.580 91.020 62.995 135.710 ;
        LAYER M3 ;
        RECT  0.600 247.660 23.220 248.740 ;
        RECT  0.600 247.660 22.900 249.400 ;
        RECT  26.260 247.660 64.400 248.740 ;
        RECT  26.580 247.660 27.000 249.400 ;
        RECT  30.440 247.660 64.400 249.400 ;
        RECT  0.600 124.090 64.400 129.850 ;
        RECT  1.640 124.090 63.600 135.790 ;
        RECT  1.810 124.090 2.830 154.520 ;
        RECT  3.510 124.090 63.600 171.560 ;
        RECT  4.040 123.970 60.900 171.560 ;
        RECT  1.640 155.040 63.600 171.560 ;
        RECT  1.640 183.580 63.600 185.950 ;
        RECT  5.515 124.090 63.600 200.820 ;
        RECT  1.640 196.170 63.600 200.820 ;
        RECT  0.600 0.600 64.400 60.480 ;
        RECT  2.000 0.000 63.000 88.700 ;
        RECT  0.600 0.600 1.480 91.220 ;
        RECT  0.600 90.750 64.400 91.220 ;
        LAYER TOP_M ;
        RECT  0.600 247.690 64.400 248.850 ;
        RECT  0.600 247.690 23.010 249.400 ;
        RECT  26.470 247.690 27.110 249.400 ;
        RECT  30.330 247.690 64.400 249.400 ;
        RECT  2.000 0.000 63.000 91.190 ;
        RECT  0.600 0.600 64.400 91.190 ;
    END
END pc3t05u

MACRO pc3t05d
    CLASS PAD ;
    FOREIGN pc3t05d 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 65.000 BY 250.000 ;
    SYMMETRY X Y R90 ;
    SITE IOSite_c ;
    PIN PAD
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 55.440  LAYER TOP_M  ;
        ANTENNAPARTIALMETALSIDEAREA 287.938  LAYER M3  ;
        ANTENNAPARTIALMETALSIDEAREA 480.740  LAYER M2  ;
        ANTENNADIFFAREA 2657.280  LAYER TOP_M  ;
        ANTENNADIFFAREA 2657.280  LAYER M3  ;
        ANTENNADIFFAREA 1209.600  LAYER M2  ;
        ANTENNAPARTIALCUTAREA 632.318  LAYER TOP_V  ;
        ANTENNAPARTIALCUTAREA 349.898  LAYER V3  ;
        ANTENNAPARTIALCUTAREA 255.798  LAYER V2  ;
        PORT
        LAYER M3 ;
        RECT  23.740 249.580 25.740 250.000 ;
        LAYER M2 ;
        RECT  2.000 61.000 63.000 90.230 ;
        RECT  23.740 246.275 25.740 250.000 ;
        END
    END PAD
    PIN OEN
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 81.726  LAYER M2  ;
        ANTENNAPARTIALMETALSIDEAREA 67.374  LAYER M1  ;
        ANTENNAPARTIALMETALSIDEAREA 41.679  LAYER M3  ;
        ANTENNADIFFAREA 0.250  LAYER M3  ;
        ANTENNAPARTIALCUTAREA 0.135  LAYER V3  ;
        ANTENNAPARTIALCUTAREA 0.203  LAYER V2  ;
        ANTENNAGATEAREA 8.100  LAYER M2  ;
        ANTENNAGATEAREA 9.900  LAYER M3  ;
        PORT
        LAYER M3 ;
        RECT  28.870 249.580 29.600 250.000 ;
        LAYER M2 ;
        RECT  28.870 249.580 29.600 250.000 ;
        END
    END OEN
    PIN I
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 67.374  LAYER M1  ;
        ANTENNAPARTIALMETALSIDEAREA 80.804  LAYER M2  ;
        ANTENNAPARTIALMETALSIDEAREA 41.096  LAYER M3  ;
        ANTENNADIFFAREA 0.250  LAYER M3  ;
        ANTENNAPARTIALCUTAREA 0.270  LAYER V2  ;
        ANTENNAPARTIALCUTAREA 0.135  LAYER V3  ;
        ANTENNAGATEAREA 18.900  LAYER M2  ;
        ANTENNAGATEAREA 20.700  LAYER M3  ;
        PORT
        LAYER M3 ;
        RECT  27.840 249.580 28.570 250.000 ;
        LAYER M2 ;
        RECT  27.840 249.580 28.570 250.000 ;
        END
    END I
    PIN VDDO
        DIRECTION INOUT ;
        USE power ;
        PORT
        LAYER M3 ;
        RECT  64.200 192.330 65.000 200.640 ;
        RECT  0.000 201.660 65.000 221.520 ;
        RECT  0.000 222.720 65.000 246.820 ;
        RECT  0.000 192.330 0.800 200.640 ;
        LAYER M2 ;
        RECT  0.000 186.470 65.000 195.650 ;
        LAYER TOP_M ;
        RECT  0.000 195.170 65.000 200.640 ;
        RECT  0.000 201.660 65.000 221.520 ;
        RECT  0.000 222.720 65.000 246.820 ;
        END
    END VDDO
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        PORT
        LAYER M3 ;
        RECT  64.200 163.510 65.000 190.890 ;
        RECT  0.000 163.510 0.800 190.890 ;
        LAYER M2 ;
        RECT  0.000 172.080 65.000 183.060 ;
        LAYER TOP_M ;
        RECT  0.000 163.500 65.000 194.560 ;
        END
    END VDD
    PIN VSSO
        DIRECTION INOUT ;
        USE ground ;
        PORT
        LAYER M3 ;
        RECT  0.000 92.060 65.000 123.250 ;
        RECT  64.200 149.940 65.000 162.610 ;
        RECT  0.000 149.940 0.800 162.610 ;
        LAYER M2 ;
        RECT  0.000 147.040 65.000 154.520 ;
        LAYER TOP_M ;
        RECT  0.000 92.060 65.000 123.250 ;
        RECT  0.000 155.410 65.000 162.610 ;
        END
    END VSSO
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        PORT
        LAYER M3 ;
        RECT  64.200 130.690 65.000 148.880 ;
        RECT  0.000 130.690 0.800 148.880 ;
        LAYER M2 ;
        RECT  0.000 136.310 65.000 146.340 ;
        LAYER TOP_M ;
        RECT  0.000 123.850 65.000 154.560 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  2.000 0.000 63.000 250.000 ;
        RECT  0.000 88.990 65.000 130.360 ;
        RECT  0.000 136.510 65.000 157.550 ;
        RECT  0.315 158.150 64.700 158.460 ;
        RECT  0.300 158.930 64.700 159.230 ;
        RECT  0.300 159.530 64.700 159.830 ;
        RECT  0.300 160.130 64.700 160.430 ;
        RECT  0.300 160.730 64.700 161.030 ;
        RECT  0.300 161.330 64.700 161.630 ;
        RECT  0.300 161.910 64.700 162.190 ;
        RECT  0.300 162.490 64.700 162.770 ;
        RECT  0.300 163.070 64.700 163.350 ;
        RECT  0.300 163.650 64.700 163.950 ;
        RECT  0.300 164.250 64.700 164.550 ;
        RECT  0.300 164.850 64.700 165.150 ;
        RECT  0.300 165.450 64.700 165.750 ;
        RECT  0.300 166.050 64.700 166.350 ;
        RECT  0.300 166.650 64.700 166.960 ;
        RECT  0.300 167.260 64.700 167.560 ;
        RECT  0.300 167.860 64.700 168.160 ;
        RECT  0.000 169.150 65.000 197.240 ;
        RECT  0.600 0.600 64.400 250.000 ;
        RECT  0.000 198.470 65.000 250.000 ;
        LAYER M2 ;
        RECT  63.180 196.430 63.670 249.400 ;
        RECT  0.600 196.440 64.400 245.485 ;
        RECT  26.530 196.440 64.400 248.790 ;
        RECT  0.600 196.440 22.950 249.400 ;
        RECT  26.530 196.440 27.050 249.400 ;
        RECT  30.390 196.440 64.400 249.400 ;
        RECT  0.600 183.850 64.400 185.680 ;
        RECT  46.230 183.850 51.730 185.870 ;
        RECT  4.480 154.920 7.530 171.290 ;
        RECT  8.170 155.125 8.490 171.290 ;
        RECT  21.210 155.160 21.560 171.290 ;
        RECT  21.860 155.140 22.180 171.290 ;
        RECT  31.895 155.120 35.765 171.290 ;
        RECT  49.255 155.125 51.495 171.290 ;
        RECT  52.435 155.295 52.745 171.290 ;
        RECT  53.655 155.035 53.935 171.290 ;
        RECT  56.365 155.280 56.645 171.290 ;
        RECT  57.120 155.300 57.400 171.290 ;
        RECT  57.835 155.130 58.115 171.290 ;
        RECT  0.600 155.310 64.400 171.290 ;
        RECT  53.895 155.310 55.870 171.370 ;
        RECT  3.170 155.310 3.450 171.380 ;
        RECT  34.655 155.310 38.715 171.480 ;
        RECT  39.605 155.310 42.020 171.480 ;
        RECT  2.000 0.000 63.000 60.210 ;
        RECT  0.600 0.600 64.400 60.210 ;
        RECT  0.600 0.600 1.210 135.520 ;
        RECT  0.600 91.020 64.400 135.520 ;
        RECT  4.080 91.020 60.940 135.690 ;
        RECT  62.580 91.020 62.995 135.710 ;
        LAYER M3 ;
        RECT  0.600 247.660 23.220 248.740 ;
        RECT  0.600 247.660 22.900 249.400 ;
        RECT  26.260 247.660 64.400 248.740 ;
        RECT  26.580 247.660 27.000 249.400 ;
        RECT  30.440 247.660 64.400 249.400 ;
        RECT  0.600 124.090 64.400 129.850 ;
        RECT  1.640 124.090 63.600 135.790 ;
        RECT  1.810 124.090 2.830 154.520 ;
        RECT  3.510 124.090 63.600 171.560 ;
        RECT  4.040 123.970 60.900 171.560 ;
        RECT  1.640 155.040 63.600 171.560 ;
        RECT  1.640 183.580 63.600 185.950 ;
        RECT  5.515 124.090 63.600 200.820 ;
        RECT  1.640 196.170 63.600 200.820 ;
        RECT  0.600 0.600 64.400 60.480 ;
        RECT  2.000 0.000 63.000 88.700 ;
        RECT  0.600 0.600 1.480 91.220 ;
        RECT  0.600 90.750 64.400 91.220 ;
        LAYER TOP_M ;
        RECT  0.600 247.690 64.400 248.850 ;
        RECT  0.600 247.690 23.010 249.400 ;
        RECT  26.470 247.690 27.110 249.400 ;
        RECT  30.330 247.690 64.400 249.400 ;
        RECT  2.000 0.000 63.000 91.190 ;
        RECT  0.600 0.600 64.400 91.190 ;
    END
END pc3t05d

MACRO pc3t05
    CLASS PAD ;
    FOREIGN pc3t05 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 65.000 BY 250.000 ;
    SYMMETRY X Y R90 ;
    SITE IOSite_c ;
    PIN PAD
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 55.440  LAYER TOP_M  ;
        ANTENNAPARTIALMETALSIDEAREA 287.938  LAYER M3  ;
        ANTENNAPARTIALMETALSIDEAREA 480.740  LAYER M2  ;
        ANTENNADIFFAREA 2657.280  LAYER TOP_M  ;
        ANTENNADIFFAREA 2657.280  LAYER M3  ;
        ANTENNADIFFAREA 1209.600  LAYER M2  ;
        ANTENNAPARTIALCUTAREA 632.318  LAYER TOP_V  ;
        ANTENNAPARTIALCUTAREA 349.898  LAYER V3  ;
        ANTENNAPARTIALCUTAREA 255.798  LAYER V2  ;
        PORT
        LAYER M3 ;
        RECT  23.740 249.580 25.740 250.000 ;
        LAYER M2 ;
        RECT  2.000 61.000 63.000 90.230 ;
        RECT  23.740 246.275 25.740 250.000 ;
        END
    END PAD
    PIN OEN
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 81.726  LAYER M2  ;
        ANTENNAPARTIALMETALSIDEAREA 67.374  LAYER M1  ;
        ANTENNAPARTIALMETALSIDEAREA 41.679  LAYER M3  ;
        ANTENNADIFFAREA 0.250  LAYER M3  ;
        ANTENNAPARTIALCUTAREA 0.203  LAYER V2  ;
        ANTENNAPARTIALCUTAREA 0.135  LAYER V3  ;
        ANTENNAGATEAREA 8.100  LAYER M2  ;
        ANTENNAGATEAREA 9.900  LAYER M3  ;
        PORT
        LAYER M3 ;
        RECT  28.870 249.580 29.600 250.000 ;
        LAYER M2 ;
        RECT  28.870 249.580 29.600 250.000 ;
        END
    END OEN
    PIN I
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 80.804  LAYER M2  ;
        ANTENNAPARTIALMETALSIDEAREA 67.374  LAYER M1  ;
        ANTENNAPARTIALMETALSIDEAREA 41.096  LAYER M3  ;
        ANTENNADIFFAREA 0.250  LAYER M3  ;
        ANTENNAPARTIALCUTAREA 0.135  LAYER V3  ;
        ANTENNAPARTIALCUTAREA 0.270  LAYER V2  ;
        ANTENNAGATEAREA 18.900  LAYER M2  ;
        ANTENNAGATEAREA 20.700  LAYER M3  ;
        PORT
        LAYER M3 ;
        RECT  27.840 249.580 28.570 250.000 ;
        LAYER M2 ;
        RECT  27.840 249.580 28.570 250.000 ;
        END
    END I
    PIN VDDO
        DIRECTION INOUT ;
        USE power ;
        PORT
        LAYER M3 ;
        RECT  64.200 192.330 65.000 200.640 ;
        RECT  0.000 201.660 65.000 221.520 ;
        RECT  0.000 222.720 65.000 246.820 ;
        RECT  0.000 192.330 0.800 200.640 ;
        LAYER M2 ;
        RECT  0.000 186.470 65.000 195.650 ;
        LAYER TOP_M ;
        RECT  0.000 195.170 65.000 200.640 ;
        RECT  0.000 201.660 65.000 221.520 ;
        RECT  0.000 222.720 65.000 246.820 ;
        END
    END VDDO
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        PORT
        LAYER M3 ;
        RECT  64.200 163.510 65.000 190.890 ;
        RECT  0.000 163.510 0.800 190.890 ;
        LAYER M2 ;
        RECT  0.000 172.080 65.000 183.060 ;
        LAYER TOP_M ;
        RECT  0.000 163.500 65.000 194.560 ;
        END
    END VDD
    PIN VSSO
        DIRECTION INOUT ;
        USE ground ;
        PORT
        LAYER M3 ;
        RECT  0.000 92.060 65.000 123.250 ;
        RECT  64.200 149.940 65.000 162.610 ;
        RECT  0.000 149.940 0.800 162.610 ;
        LAYER M2 ;
        RECT  0.000 147.040 65.000 154.520 ;
        LAYER TOP_M ;
        RECT  0.000 92.060 65.000 123.250 ;
        RECT  0.000 155.410 65.000 162.610 ;
        END
    END VSSO
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        PORT
        LAYER M3 ;
        RECT  64.200 130.690 65.000 148.880 ;
        RECT  0.000 130.690 0.800 148.880 ;
        LAYER M2 ;
        RECT  0.000 136.310 65.000 146.340 ;
        LAYER TOP_M ;
        RECT  0.000 123.850 65.000 154.560 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  2.000 0.000 63.000 250.000 ;
        RECT  0.000 88.990 65.000 130.360 ;
        RECT  0.000 136.510 65.000 157.550 ;
        RECT  0.315 158.150 64.700 158.460 ;
        RECT  0.300 158.930 64.700 159.230 ;
        RECT  0.300 159.530 64.700 159.830 ;
        RECT  0.300 160.130 64.700 160.430 ;
        RECT  0.300 160.730 64.700 161.030 ;
        RECT  0.300 161.330 64.700 161.630 ;
        RECT  0.300 161.910 64.700 162.190 ;
        RECT  0.300 162.490 64.700 162.770 ;
        RECT  0.300 163.070 64.700 163.350 ;
        RECT  0.300 163.650 64.700 163.950 ;
        RECT  0.300 164.250 64.700 164.550 ;
        RECT  0.300 164.850 64.700 165.150 ;
        RECT  0.300 165.450 64.700 165.750 ;
        RECT  0.300 166.050 64.700 166.350 ;
        RECT  0.300 166.650 64.700 166.960 ;
        RECT  0.300 167.260 64.700 167.560 ;
        RECT  0.300 167.860 64.700 168.160 ;
        RECT  0.000 169.150 65.000 197.240 ;
        RECT  0.600 0.600 64.400 250.000 ;
        RECT  0.000 198.470 65.000 250.000 ;
        LAYER M2 ;
        RECT  63.180 196.430 63.670 249.400 ;
        RECT  0.600 196.440 64.400 245.485 ;
        RECT  26.530 196.440 64.400 248.790 ;
        RECT  0.600 196.440 22.950 249.400 ;
        RECT  26.530 196.440 27.050 249.400 ;
        RECT  30.390 196.440 64.400 249.400 ;
        RECT  0.600 183.850 64.400 185.680 ;
        RECT  46.230 183.850 51.730 185.870 ;
        RECT  4.480 154.920 7.530 171.290 ;
        RECT  8.170 155.125 8.490 171.290 ;
        RECT  21.210 155.160 21.560 171.290 ;
        RECT  21.860 155.140 22.180 171.290 ;
        RECT  31.895 155.120 35.765 171.290 ;
        RECT  53.655 155.035 53.935 171.290 ;
        RECT  56.365 155.280 56.645 171.290 ;
        RECT  57.120 155.300 57.400 171.290 ;
        RECT  57.835 155.130 58.115 171.290 ;
        RECT  0.600 155.310 64.400 171.290 ;
        RECT  53.895 155.310 55.870 171.370 ;
        RECT  3.170 155.310 3.450 171.380 ;
        RECT  34.655 155.310 38.715 171.480 ;
        RECT  39.605 155.310 42.020 171.480 ;
        RECT  2.000 0.000 63.000 60.210 ;
        RECT  0.600 0.600 64.400 60.210 ;
        RECT  0.600 0.600 1.210 135.520 ;
        RECT  0.600 91.020 64.400 135.520 ;
        RECT  4.080 91.020 60.940 135.690 ;
        RECT  62.580 91.020 62.995 135.710 ;
        LAYER M3 ;
        RECT  0.600 247.660 23.220 248.740 ;
        RECT  0.600 247.660 22.900 249.400 ;
        RECT  26.260 247.660 64.400 248.740 ;
        RECT  26.580 247.660 27.000 249.400 ;
        RECT  30.440 247.660 64.400 249.400 ;
        RECT  0.600 124.090 64.400 129.850 ;
        RECT  1.640 124.090 63.600 135.790 ;
        RECT  1.810 124.090 2.830 154.520 ;
        RECT  3.510 124.090 63.600 171.560 ;
        RECT  4.040 123.970 60.900 171.560 ;
        RECT  1.640 155.040 63.600 171.560 ;
        RECT  1.640 183.580 63.600 185.950 ;
        RECT  5.515 124.090 63.600 200.820 ;
        RECT  1.640 196.170 63.600 200.820 ;
        RECT  0.600 0.600 64.400 60.480 ;
        RECT  2.000 0.000 63.000 88.700 ;
        RECT  0.600 0.600 1.480 91.220 ;
        RECT  0.600 90.750 64.400 91.220 ;
        LAYER TOP_M ;
        RECT  0.600 247.690 64.400 248.850 ;
        RECT  0.600 247.690 23.010 249.400 ;
        RECT  26.470 247.690 27.110 249.400 ;
        RECT  30.330 247.690 64.400 249.400 ;
        RECT  2.000 0.000 63.000 91.190 ;
        RECT  0.600 0.600 64.400 91.190 ;
    END
END pc3t05

MACRO pc3t04u
    CLASS PAD ;
    FOREIGN pc3t04u 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 65.000 BY 250.000 ;
    SYMMETRY X Y R90 ;
    SITE IOSite_c ;
    PIN PAD
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 55.440  LAYER TOP_M  ;
        ANTENNAPARTIALMETALSIDEAREA 287.938  LAYER M3  ;
        ANTENNAPARTIALMETALSIDEAREA 480.740  LAYER M2  ;
        ANTENNADIFFAREA 2657.280  LAYER TOP_M  ;
        ANTENNADIFFAREA 2657.280  LAYER M3  ;
        ANTENNADIFFAREA 1209.600  LAYER M2  ;
        ANTENNAPARTIALCUTAREA 632.318  LAYER TOP_V  ;
        ANTENNAPARTIALCUTAREA 349.898  LAYER V3  ;
        ANTENNAPARTIALCUTAREA 255.798  LAYER V2  ;
        PORT
        LAYER M3 ;
        RECT  23.740 249.580 25.740 250.000 ;
        LAYER M2 ;
        RECT  2.000 61.000 63.000 90.230 ;
        RECT  23.740 246.275 25.740 250.000 ;
        END
    END PAD
    PIN OEN
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 81.726  LAYER M2  ;
        ANTENNAPARTIALMETALSIDEAREA 67.374  LAYER M1  ;
        ANTENNAPARTIALMETALSIDEAREA 41.679  LAYER M3  ;
        ANTENNADIFFAREA 0.250  LAYER M3  ;
        ANTENNAPARTIALCUTAREA 0.203  LAYER V2  ;
        ANTENNAPARTIALCUTAREA 0.135  LAYER V3  ;
        ANTENNAGATEAREA 8.100  LAYER M2  ;
        ANTENNAGATEAREA 9.900  LAYER M3  ;
        PORT
        LAYER M3 ;
        RECT  28.870 249.580 29.600 250.000 ;
        LAYER M2 ;
        RECT  28.870 249.580 29.600 250.000 ;
        END
    END OEN
    PIN I
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 67.374  LAYER M1  ;
        ANTENNAPARTIALMETALSIDEAREA 80.804  LAYER M2  ;
        ANTENNAPARTIALMETALSIDEAREA 41.096  LAYER M3  ;
        ANTENNADIFFAREA 0.250  LAYER M3  ;
        ANTENNAPARTIALCUTAREA 0.270  LAYER V2  ;
        ANTENNAPARTIALCUTAREA 0.135  LAYER V3  ;
        ANTENNAGATEAREA 18.900  LAYER M2  ;
        ANTENNAGATEAREA 20.700  LAYER M3  ;
        PORT
        LAYER M3 ;
        RECT  27.840 249.580 28.570 250.000 ;
        LAYER M2 ;
        RECT  27.840 249.580 28.570 250.000 ;
        END
    END I
    PIN VDDO
        DIRECTION INOUT ;
        USE power ;
        PORT
        LAYER M3 ;
        RECT  64.200 192.330 65.000 200.640 ;
        RECT  0.000 201.660 65.000 221.520 ;
        RECT  0.000 222.720 65.000 246.820 ;
        RECT  0.000 192.330 0.800 200.640 ;
        LAYER M2 ;
        RECT  0.000 186.470 65.000 195.650 ;
        LAYER TOP_M ;
        RECT  0.000 195.170 65.000 200.640 ;
        RECT  0.000 201.660 65.000 221.520 ;
        RECT  0.000 222.720 65.000 246.820 ;
        END
    END VDDO
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        PORT
        LAYER M3 ;
        RECT  64.200 163.510 65.000 190.890 ;
        RECT  0.000 163.510 0.800 190.890 ;
        LAYER M2 ;
        RECT  0.000 172.080 65.000 183.060 ;
        LAYER TOP_M ;
        RECT  0.000 163.500 65.000 194.560 ;
        END
    END VDD
    PIN VSSO
        DIRECTION INOUT ;
        USE ground ;
        PORT
        LAYER M3 ;
        RECT  0.000 92.060 65.000 123.250 ;
        RECT  64.200 149.940 65.000 162.610 ;
        RECT  0.000 149.940 0.800 162.610 ;
        LAYER M2 ;
        RECT  0.000 147.040 65.000 154.520 ;
        LAYER TOP_M ;
        RECT  0.000 92.060 65.000 123.250 ;
        RECT  0.000 155.410 65.000 162.610 ;
        END
    END VSSO
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        PORT
        LAYER M3 ;
        RECT  64.200 130.690 65.000 148.880 ;
        RECT  0.000 130.690 0.800 148.880 ;
        LAYER M2 ;
        RECT  0.000 136.310 65.000 146.340 ;
        LAYER TOP_M ;
        RECT  0.000 123.850 65.000 154.560 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  2.000 0.000 63.000 250.000 ;
        RECT  0.000 88.990 65.000 130.360 ;
        RECT  0.000 136.510 65.000 157.550 ;
        RECT  0.315 158.150 64.700 158.460 ;
        RECT  0.300 158.930 64.700 159.230 ;
        RECT  0.300 159.530 64.700 159.830 ;
        RECT  0.300 160.130 64.700 160.430 ;
        RECT  0.300 160.730 64.700 161.030 ;
        RECT  0.300 161.330 64.700 161.630 ;
        RECT  0.300 161.910 64.700 162.190 ;
        RECT  0.300 162.490 64.700 162.770 ;
        RECT  0.300 163.070 64.700 163.350 ;
        RECT  0.300 163.650 64.700 163.950 ;
        RECT  0.300 164.250 64.700 164.550 ;
        RECT  0.300 164.850 64.700 165.150 ;
        RECT  0.300 165.450 64.700 165.750 ;
        RECT  0.300 166.050 64.700 166.350 ;
        RECT  0.300 166.650 64.700 166.960 ;
        RECT  0.300 167.260 64.700 167.560 ;
        RECT  0.300 167.860 64.700 168.160 ;
        RECT  0.000 169.150 65.000 197.240 ;
        RECT  0.600 0.600 64.400 250.000 ;
        RECT  0.000 198.470 65.000 250.000 ;
        LAYER M2 ;
        RECT  63.180 196.430 63.670 249.400 ;
        RECT  0.600 196.440 64.400 245.485 ;
        RECT  26.530 196.440 64.400 248.790 ;
        RECT  0.600 196.440 22.950 249.400 ;
        RECT  26.530 196.440 27.050 249.400 ;
        RECT  30.390 196.440 64.400 249.400 ;
        RECT  0.600 183.850 64.400 185.680 ;
        RECT  46.230 183.850 51.730 185.870 ;
        RECT  4.830 155.120 7.380 171.290 ;
        RECT  8.170 155.125 8.490 171.290 ;
        RECT  21.140 155.160 21.490 171.290 ;
        RECT  21.790 155.140 22.110 171.290 ;
        RECT  53.655 155.035 53.935 171.290 ;
        RECT  56.365 155.280 56.645 171.290 ;
        RECT  57.120 155.300 57.400 171.290 ;
        RECT  57.835 155.130 58.115 171.290 ;
        RECT  0.600 155.310 64.400 171.290 ;
        RECT  53.895 155.310 55.870 171.370 ;
        RECT  33.280 155.310 33.780 171.375 ;
        RECT  3.170 155.310 3.450 171.380 ;
        RECT  34.655 155.310 38.715 171.480 ;
        RECT  39.605 155.310 42.020 171.480 ;
        RECT  2.000 0.000 63.000 60.210 ;
        RECT  0.600 0.600 64.400 60.210 ;
        RECT  0.600 0.600 1.210 135.520 ;
        RECT  0.600 91.020 64.400 135.520 ;
        RECT  4.080 91.020 60.940 135.690 ;
        RECT  62.580 91.020 62.995 135.710 ;
        LAYER M3 ;
        RECT  0.600 247.660 23.220 248.740 ;
        RECT  0.600 247.660 22.900 249.400 ;
        RECT  26.260 247.660 64.400 248.740 ;
        RECT  26.580 247.660 27.000 249.400 ;
        RECT  30.440 247.660 64.400 249.400 ;
        RECT  0.600 124.090 64.400 129.850 ;
        RECT  1.640 124.090 63.600 135.790 ;
        RECT  1.810 124.090 2.830 154.520 ;
        RECT  3.195 124.090 63.600 171.560 ;
        RECT  3.325 123.900 61.330 171.560 ;
        RECT  1.640 155.040 63.600 171.560 ;
        RECT  1.640 183.580 63.600 185.950 ;
        RECT  5.515 124.090 63.600 200.820 ;
        RECT  1.640 196.170 63.600 200.820 ;
        RECT  0.600 0.600 64.400 60.480 ;
        RECT  2.000 0.000 63.000 88.700 ;
        RECT  0.600 0.600 1.480 91.220 ;
        RECT  0.600 90.750 64.400 91.220 ;
        LAYER TOP_M ;
        RECT  0.600 247.690 64.400 248.850 ;
        RECT  0.600 247.690 23.010 249.400 ;
        RECT  26.470 247.690 27.110 249.400 ;
        RECT  30.330 247.690 64.400 249.400 ;
        RECT  2.000 0.000 63.000 91.190 ;
        RECT  0.600 0.600 64.400 91.190 ;
    END
END pc3t04u

MACRO pc3t04d
    CLASS PAD ;
    FOREIGN pc3t04d 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 65.000 BY 250.000 ;
    SYMMETRY X Y R90 ;
    SITE IOSite_c ;
    PIN PAD
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 55.440  LAYER TOP_M  ;
        ANTENNAPARTIALMETALSIDEAREA 287.938  LAYER M3  ;
        ANTENNAPARTIALMETALSIDEAREA 480.740  LAYER M2  ;
        ANTENNADIFFAREA 2657.280  LAYER TOP_M  ;
        ANTENNADIFFAREA 2657.280  LAYER M3  ;
        ANTENNADIFFAREA 1209.600  LAYER M2  ;
        ANTENNAPARTIALCUTAREA 632.318  LAYER TOP_V  ;
        ANTENNAPARTIALCUTAREA 349.898  LAYER V3  ;
        ANTENNAPARTIALCUTAREA 255.798  LAYER V2  ;
        PORT
        LAYER M3 ;
        RECT  23.740 249.580 25.740 250.000 ;
        LAYER M2 ;
        RECT  2.000 61.000 63.000 90.230 ;
        RECT  23.740 246.275 25.740 250.000 ;
        END
    END PAD
    PIN OEN
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 81.726  LAYER M2  ;
        ANTENNAPARTIALMETALSIDEAREA 67.374  LAYER M1  ;
        ANTENNAPARTIALMETALSIDEAREA 41.679  LAYER M3  ;
        ANTENNADIFFAREA 0.250  LAYER M3  ;
        ANTENNAPARTIALCUTAREA 0.203  LAYER V2  ;
        ANTENNAPARTIALCUTAREA 0.135  LAYER V3  ;
        ANTENNAGATEAREA 8.100  LAYER M2  ;
        ANTENNAGATEAREA 9.900  LAYER M3  ;
        PORT
        LAYER M3 ;
        RECT  28.870 249.580 29.600 250.000 ;
        LAYER M2 ;
        RECT  28.870 249.580 29.600 250.000 ;
        END
    END OEN
    PIN I
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 67.374  LAYER M1  ;
        ANTENNAPARTIALMETALSIDEAREA 80.804  LAYER M2  ;
        ANTENNAPARTIALMETALSIDEAREA 41.096  LAYER M3  ;
        ANTENNADIFFAREA 0.250  LAYER M3  ;
        ANTENNAPARTIALCUTAREA 0.270  LAYER V2  ;
        ANTENNAPARTIALCUTAREA 0.135  LAYER V3  ;
        ANTENNAGATEAREA 18.900  LAYER M2  ;
        ANTENNAGATEAREA 20.700  LAYER M3  ;
        PORT
        LAYER M3 ;
        RECT  27.840 249.580 28.570 250.000 ;
        LAYER M2 ;
        RECT  27.840 249.580 28.570 250.000 ;
        END
    END I
    PIN VDDO
        DIRECTION INOUT ;
        USE power ;
        PORT
        LAYER M3 ;
        RECT  64.200 192.330 65.000 200.640 ;
        RECT  0.000 201.660 65.000 221.520 ;
        RECT  0.000 222.720 65.000 246.820 ;
        RECT  0.000 192.330 0.800 200.640 ;
        LAYER M2 ;
        RECT  0.000 186.470 65.000 195.650 ;
        LAYER TOP_M ;
        RECT  0.000 195.170 65.000 200.640 ;
        RECT  0.000 201.660 65.000 221.520 ;
        RECT  0.000 222.720 65.000 246.820 ;
        END
    END VDDO
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        PORT
        LAYER M3 ;
        RECT  64.200 163.510 65.000 190.890 ;
        RECT  0.000 163.510 0.800 190.890 ;
        LAYER M2 ;
        RECT  0.000 172.080 65.000 183.060 ;
        LAYER TOP_M ;
        RECT  0.000 163.500 65.000 194.560 ;
        END
    END VDD
    PIN VSSO
        DIRECTION INOUT ;
        USE ground ;
        PORT
        LAYER M3 ;
        RECT  0.000 92.060 65.000 123.250 ;
        RECT  64.200 149.940 65.000 162.610 ;
        RECT  0.000 149.940 0.800 162.610 ;
        LAYER M2 ;
        RECT  0.000 147.040 65.000 154.520 ;
        LAYER TOP_M ;
        RECT  0.000 92.060 65.000 123.250 ;
        RECT  0.000 155.410 65.000 162.610 ;
        END
    END VSSO
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        PORT
        LAYER M3 ;
        RECT  64.200 130.690 65.000 148.880 ;
        RECT  0.000 130.690 0.800 148.880 ;
        LAYER M2 ;
        RECT  0.000 136.310 65.000 146.340 ;
        LAYER TOP_M ;
        RECT  0.000 123.850 65.000 154.560 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  2.000 0.000 63.000 250.000 ;
        RECT  0.000 88.990 65.000 130.360 ;
        RECT  0.000 136.510 65.000 157.550 ;
        RECT  0.315 158.150 64.700 158.460 ;
        RECT  0.300 158.930 64.700 159.230 ;
        RECT  0.300 159.530 64.700 159.830 ;
        RECT  0.300 160.130 64.700 160.430 ;
        RECT  0.300 160.730 64.700 161.030 ;
        RECT  0.300 161.330 64.700 161.630 ;
        RECT  0.300 161.910 64.700 162.190 ;
        RECT  0.300 162.490 64.700 162.770 ;
        RECT  0.300 163.070 64.700 163.350 ;
        RECT  0.300 163.650 64.700 163.950 ;
        RECT  0.300 164.250 64.700 164.550 ;
        RECT  0.300 164.850 64.700 165.150 ;
        RECT  0.300 165.450 64.700 165.750 ;
        RECT  0.300 166.050 64.700 166.350 ;
        RECT  0.300 166.650 64.700 166.960 ;
        RECT  0.300 167.260 64.700 167.560 ;
        RECT  0.300 167.860 64.700 168.160 ;
        RECT  0.000 169.150 65.000 197.240 ;
        RECT  0.600 0.600 64.400 250.000 ;
        RECT  0.000 198.470 65.000 250.000 ;
        LAYER M2 ;
        RECT  63.180 196.430 63.670 249.400 ;
        RECT  0.600 196.440 64.400 245.485 ;
        RECT  26.530 196.440 64.400 248.790 ;
        RECT  0.600 196.440 22.950 249.400 ;
        RECT  26.530 196.440 27.050 249.400 ;
        RECT  30.390 196.440 64.400 249.400 ;
        RECT  0.600 183.850 64.400 185.680 ;
        RECT  46.230 183.850 51.730 185.870 ;
        RECT  4.830 155.120 7.380 171.290 ;
        RECT  8.170 155.125 8.490 171.290 ;
        RECT  21.140 155.160 21.490 171.290 ;
        RECT  21.790 155.140 22.110 171.290 ;
        RECT  49.425 155.125 51.665 171.290 ;
        RECT  52.605 155.295 52.915 171.290 ;
        RECT  53.655 155.035 53.935 171.290 ;
        RECT  56.365 155.280 56.645 171.290 ;
        RECT  57.120 155.300 57.400 171.290 ;
        RECT  57.835 155.130 58.115 171.290 ;
        RECT  0.600 155.310 64.400 171.290 ;
        RECT  53.895 155.310 55.870 171.370 ;
        RECT  3.170 155.310 3.450 171.380 ;
        RECT  34.655 155.310 38.715 171.480 ;
        RECT  39.605 155.310 42.020 171.480 ;
        RECT  2.000 0.000 63.000 60.210 ;
        RECT  0.600 0.600 64.400 60.210 ;
        RECT  0.600 0.600 1.210 135.520 ;
        RECT  0.600 91.020 64.400 135.520 ;
        RECT  4.080 91.020 60.940 135.690 ;
        RECT  62.580 91.020 62.995 135.710 ;
        LAYER M3 ;
        RECT  0.600 247.660 23.220 248.740 ;
        RECT  0.600 247.660 22.900 249.400 ;
        RECT  26.260 247.660 64.400 248.740 ;
        RECT  26.580 247.660 27.000 249.400 ;
        RECT  30.440 247.660 64.400 249.400 ;
        RECT  0.600 124.090 64.400 129.850 ;
        RECT  1.640 124.090 63.600 135.790 ;
        RECT  1.810 124.090 2.830 154.520 ;
        RECT  3.195 124.090 63.600 171.560 ;
        RECT  3.325 123.900 61.330 171.560 ;
        RECT  1.640 155.040 63.600 171.560 ;
        RECT  1.640 183.580 63.600 185.950 ;
        RECT  5.515 124.090 63.600 200.820 ;
        RECT  1.640 196.170 63.600 200.820 ;
        RECT  0.600 0.600 64.400 60.480 ;
        RECT  2.000 0.000 63.000 88.700 ;
        RECT  0.600 0.600 1.480 91.220 ;
        RECT  0.600 90.750 64.400 91.220 ;
        LAYER TOP_M ;
        RECT  0.600 247.690 64.400 248.850 ;
        RECT  0.600 247.690 23.010 249.400 ;
        RECT  26.470 247.690 27.110 249.400 ;
        RECT  30.330 247.690 64.400 249.400 ;
        RECT  2.000 0.000 63.000 91.190 ;
        RECT  0.600 0.600 64.400 91.190 ;
    END
END pc3t04d

MACRO pc3t04
    CLASS PAD ;
    FOREIGN pc3t04 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 65.000 BY 250.000 ;
    SYMMETRY X Y R90 ;
    SITE IOSite_c ;
    PIN PAD
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 55.440  LAYER TOP_M  ;
        ANTENNAPARTIALMETALSIDEAREA 287.938  LAYER M3  ;
        ANTENNAPARTIALMETALSIDEAREA 480.740  LAYER M2  ;
        ANTENNADIFFAREA 2657.280  LAYER TOP_M  ;
        ANTENNADIFFAREA 2657.280  LAYER M3  ;
        ANTENNADIFFAREA 1209.600  LAYER M2  ;
        ANTENNAPARTIALCUTAREA 632.318  LAYER TOP_V  ;
        ANTENNAPARTIALCUTAREA 349.898  LAYER V3  ;
        ANTENNAPARTIALCUTAREA 255.798  LAYER V2  ;
        PORT
        LAYER M3 ;
        RECT  23.740 249.580 25.740 250.000 ;
        LAYER M2 ;
        RECT  2.000 61.000 63.000 90.230 ;
        RECT  23.740 246.275 25.740 250.000 ;
        END
    END PAD
    PIN OEN
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 67.374  LAYER M1  ;
        ANTENNAPARTIALMETALSIDEAREA 81.726  LAYER M2  ;
        ANTENNAPARTIALMETALSIDEAREA 41.679  LAYER M3  ;
        ANTENNADIFFAREA 0.250  LAYER M3  ;
        ANTENNAPARTIALCUTAREA 0.203  LAYER V2  ;
        ANTENNAPARTIALCUTAREA 0.135  LAYER V3  ;
        ANTENNAGATEAREA 8.100  LAYER M2  ;
        ANTENNAGATEAREA 9.900  LAYER M3  ;
        PORT
        LAYER M3 ;
        RECT  28.870 249.580 29.600 250.000 ;
        LAYER M2 ;
        RECT  28.870 249.580 29.600 250.000 ;
        END
    END OEN
    PIN I
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 67.374  LAYER M1  ;
        ANTENNAPARTIALMETALSIDEAREA 80.804  LAYER M2  ;
        ANTENNAPARTIALMETALSIDEAREA 41.096  LAYER M3  ;
        ANTENNADIFFAREA 0.250  LAYER M3  ;
        ANTENNAPARTIALCUTAREA 0.270  LAYER V2  ;
        ANTENNAPARTIALCUTAREA 0.135  LAYER V3  ;
        ANTENNAGATEAREA 18.900  LAYER M2  ;
        ANTENNAGATEAREA 20.700  LAYER M3  ;
        PORT
        LAYER M3 ;
        RECT  27.840 249.580 28.570 250.000 ;
        LAYER M2 ;
        RECT  27.840 249.580 28.570 250.000 ;
        END
    END I
    PIN VDDO
        DIRECTION INOUT ;
        USE power ;
        PORT
        LAYER M3 ;
        RECT  64.200 192.330 65.000 200.640 ;
        RECT  0.000 201.660 65.000 221.520 ;
        RECT  0.000 222.720 65.000 246.820 ;
        RECT  0.000 192.330 0.800 200.640 ;
        LAYER M2 ;
        RECT  0.000 186.470 65.000 195.650 ;
        LAYER TOP_M ;
        RECT  0.000 195.170 65.000 200.640 ;
        RECT  0.000 201.660 65.000 221.520 ;
        RECT  0.000 222.720 65.000 246.820 ;
        END
    END VDDO
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        PORT
        LAYER M3 ;
        RECT  64.200 163.510 65.000 190.890 ;
        RECT  0.000 163.510 0.800 190.890 ;
        LAYER M2 ;
        RECT  0.000 172.080 65.000 183.060 ;
        LAYER TOP_M ;
        RECT  0.000 163.500 65.000 194.560 ;
        END
    END VDD
    PIN VSSO
        DIRECTION INOUT ;
        USE ground ;
        PORT
        LAYER M3 ;
        RECT  0.000 92.060 65.000 123.250 ;
        RECT  64.200 149.940 65.000 162.610 ;
        RECT  0.000 149.940 0.800 162.610 ;
        LAYER M2 ;
        RECT  0.000 147.040 65.000 154.520 ;
        LAYER TOP_M ;
        RECT  0.000 92.060 65.000 123.250 ;
        RECT  0.000 155.410 65.000 162.610 ;
        END
    END VSSO
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        PORT
        LAYER M3 ;
        RECT  64.200 130.690 65.000 148.880 ;
        RECT  0.000 130.690 0.800 148.880 ;
        LAYER M2 ;
        RECT  0.000 136.310 65.000 146.340 ;
        LAYER TOP_M ;
        RECT  0.000 123.850 65.000 154.560 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  2.000 0.000 63.000 250.000 ;
        RECT  0.000 88.990 65.000 130.360 ;
        RECT  0.000 136.510 65.000 157.550 ;
        RECT  0.315 158.150 64.700 158.460 ;
        RECT  0.300 158.930 64.700 159.230 ;
        RECT  0.300 159.530 64.700 159.830 ;
        RECT  0.300 160.130 64.700 160.430 ;
        RECT  0.300 160.730 64.700 161.030 ;
        RECT  0.300 161.330 64.700 161.630 ;
        RECT  0.300 161.910 64.700 162.190 ;
        RECT  0.300 162.490 64.700 162.770 ;
        RECT  0.300 163.070 64.700 163.350 ;
        RECT  0.300 163.650 64.700 163.950 ;
        RECT  0.300 164.250 64.700 164.550 ;
        RECT  0.300 164.850 64.700 165.150 ;
        RECT  0.300 165.450 64.700 165.750 ;
        RECT  0.300 166.050 64.700 166.350 ;
        RECT  0.300 166.650 64.700 166.960 ;
        RECT  0.300 167.260 64.700 167.560 ;
        RECT  0.300 167.860 64.700 168.160 ;
        RECT  0.000 169.150 65.000 197.240 ;
        RECT  0.600 0.600 64.400 250.000 ;
        RECT  0.000 198.470 65.000 250.000 ;
        LAYER M2 ;
        RECT  63.180 196.430 63.670 249.400 ;
        RECT  0.600 196.440 64.400 245.485 ;
        RECT  26.530 196.440 64.400 248.790 ;
        RECT  0.600 196.440 22.950 249.400 ;
        RECT  26.530 196.440 27.050 249.400 ;
        RECT  30.390 196.440 64.400 249.400 ;
        RECT  0.600 183.850 64.400 185.680 ;
        RECT  46.230 183.850 51.730 185.870 ;
        RECT  4.830 155.120 7.380 171.290 ;
        RECT  8.170 155.125 8.490 171.290 ;
        RECT  21.140 155.160 21.490 171.290 ;
        RECT  21.790 155.140 22.110 171.290 ;
        RECT  53.655 155.035 53.935 171.290 ;
        RECT  56.365 155.280 56.645 171.290 ;
        RECT  57.120 155.300 57.400 171.290 ;
        RECT  57.835 155.130 58.115 171.290 ;
        RECT  0.600 155.310 64.400 171.290 ;
        RECT  53.895 155.310 55.870 171.370 ;
        RECT  3.170 155.310 3.450 171.380 ;
        RECT  34.655 155.310 38.715 171.480 ;
        RECT  39.605 155.310 42.020 171.480 ;
        RECT  2.000 0.000 63.000 60.210 ;
        RECT  0.600 0.600 64.400 60.210 ;
        RECT  0.600 0.600 1.210 135.520 ;
        RECT  0.600 91.020 64.400 135.520 ;
        RECT  4.080 91.020 60.940 135.690 ;
        RECT  62.580 91.020 62.995 135.710 ;
        LAYER M3 ;
        RECT  0.600 247.660 23.220 248.740 ;
        RECT  0.600 247.660 22.900 249.400 ;
        RECT  26.260 247.660 64.400 248.740 ;
        RECT  26.580 247.660 27.000 249.400 ;
        RECT  30.440 247.660 64.400 249.400 ;
        RECT  0.600 124.090 64.400 129.850 ;
        RECT  1.640 124.090 63.600 135.790 ;
        RECT  1.810 124.090 2.830 154.520 ;
        RECT  3.195 124.090 63.600 171.560 ;
        RECT  3.325 123.900 61.330 171.560 ;
        RECT  1.640 155.040 63.600 171.560 ;
        RECT  1.640 183.580 63.600 185.950 ;
        RECT  5.515 124.090 63.600 200.820 ;
        RECT  1.640 196.170 63.600 200.820 ;
        RECT  0.600 0.600 64.400 60.480 ;
        RECT  2.000 0.000 63.000 88.700 ;
        RECT  0.600 0.600 1.480 91.220 ;
        RECT  0.600 90.750 64.400 91.220 ;
        LAYER TOP_M ;
        RECT  0.600 247.690 64.400 248.850 ;
        RECT  0.600 247.690 23.010 249.400 ;
        RECT  26.470 247.690 27.110 249.400 ;
        RECT  30.330 247.690 64.400 249.400 ;
        RECT  2.000 0.000 63.000 91.190 ;
        RECT  0.600 0.600 64.400 91.190 ;
    END
END pc3t04

MACRO pc3t03u
    CLASS PAD ;
    FOREIGN pc3t03u 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 65.000 BY 250.000 ;
    SYMMETRY X Y R90 ;
    SITE IOSite_c ;
    PIN PAD
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 55.440  LAYER TOP_M  ;
        ANTENNAPARTIALMETALSIDEAREA 287.938  LAYER M3  ;
        ANTENNAPARTIALMETALSIDEAREA 480.740  LAYER M2  ;
        ANTENNADIFFAREA 2657.280  LAYER TOP_M  ;
        ANTENNADIFFAREA 2657.280  LAYER M3  ;
        ANTENNADIFFAREA 1209.600  LAYER M2  ;
        ANTENNAPARTIALCUTAREA 632.318  LAYER TOP_V  ;
        ANTENNAPARTIALCUTAREA 349.898  LAYER V3  ;
        ANTENNAPARTIALCUTAREA 255.798  LAYER V2  ;
        PORT
        LAYER M3 ;
        RECT  23.740 249.580 25.740 250.000 ;
        LAYER M2 ;
        RECT  2.000 61.000 63.000 90.230 ;
        RECT  23.740 246.275 25.740 250.000 ;
        END
    END PAD
    PIN OEN
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 67.374  LAYER M1  ;
        ANTENNAPARTIALMETALSIDEAREA 81.726  LAYER M2  ;
        ANTENNAPARTIALMETALSIDEAREA 41.679  LAYER M3  ;
        ANTENNADIFFAREA 0.250  LAYER M3  ;
        ANTENNAPARTIALCUTAREA 0.203  LAYER V2  ;
        ANTENNAPARTIALCUTAREA 0.135  LAYER V3  ;
        ANTENNAGATEAREA 8.100  LAYER M2  ;
        ANTENNAGATEAREA 9.900  LAYER M3  ;
        PORT
        LAYER M3 ;
        RECT  28.870 249.580 29.600 250.000 ;
        LAYER M2 ;
        RECT  28.870 249.580 29.600 250.000 ;
        END
    END OEN
    PIN I
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 80.804  LAYER M2  ;
        ANTENNAPARTIALMETALSIDEAREA 67.374  LAYER M1  ;
        ANTENNAPARTIALMETALSIDEAREA 41.096  LAYER M3  ;
        ANTENNADIFFAREA 0.250  LAYER M3  ;
        ANTENNAPARTIALCUTAREA 0.135  LAYER V3  ;
        ANTENNAPARTIALCUTAREA 0.270  LAYER V2  ;
        ANTENNAGATEAREA 18.900  LAYER M2  ;
        ANTENNAGATEAREA 20.700  LAYER M3  ;
        PORT
        LAYER M3 ;
        RECT  27.840 249.580 28.570 250.000 ;
        LAYER M2 ;
        RECT  27.840 249.580 28.570 250.000 ;
        END
    END I
    PIN VDDO
        DIRECTION INOUT ;
        USE power ;
        PORT
        LAYER M3 ;
        RECT  64.200 192.330 65.000 200.640 ;
        RECT  0.000 201.660 65.000 221.520 ;
        RECT  0.000 222.720 65.000 246.820 ;
        RECT  0.000 192.330 0.800 200.640 ;
        LAYER M2 ;
        RECT  0.000 186.470 65.000 195.650 ;
        LAYER TOP_M ;
        RECT  0.000 195.170 65.000 200.640 ;
        RECT  0.000 201.660 65.000 221.520 ;
        RECT  0.000 222.720 65.000 246.820 ;
        END
    END VDDO
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        PORT
        LAYER M3 ;
        RECT  64.200 163.510 65.000 190.890 ;
        RECT  0.000 163.510 0.800 190.890 ;
        LAYER M2 ;
        RECT  0.000 172.080 65.000 183.060 ;
        LAYER TOP_M ;
        RECT  0.000 163.500 65.000 194.560 ;
        END
    END VDD
    PIN VSSO
        DIRECTION INOUT ;
        USE ground ;
        PORT
        LAYER M3 ;
        RECT  0.000 92.060 65.000 123.250 ;
        RECT  64.200 149.940 65.000 162.610 ;
        RECT  0.000 149.940 0.800 162.610 ;
        LAYER M2 ;
        RECT  0.000 147.040 65.000 154.520 ;
        LAYER TOP_M ;
        RECT  0.000 92.060 65.000 123.250 ;
        RECT  0.000 155.410 65.000 162.610 ;
        END
    END VSSO
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        PORT
        LAYER M3 ;
        RECT  64.200 130.690 65.000 148.880 ;
        RECT  0.000 130.690 0.800 148.880 ;
        LAYER M2 ;
        RECT  0.000 136.310 65.000 146.340 ;
        LAYER TOP_M ;
        RECT  0.000 123.850 65.000 154.560 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  2.000 0.000 63.000 250.000 ;
        RECT  0.000 88.990 65.000 130.360 ;
        RECT  0.000 136.510 65.000 157.550 ;
        RECT  0.315 158.150 64.700 158.460 ;
        RECT  0.300 158.930 64.700 159.230 ;
        RECT  0.300 159.530 64.700 159.830 ;
        RECT  0.300 160.130 64.700 160.430 ;
        RECT  0.300 160.730 64.700 161.030 ;
        RECT  0.300 161.330 64.700 161.630 ;
        RECT  0.300 161.910 64.700 162.190 ;
        RECT  0.300 162.490 64.700 162.770 ;
        RECT  0.300 163.070 64.700 163.350 ;
        RECT  0.300 163.650 64.700 163.950 ;
        RECT  0.300 164.250 64.700 164.550 ;
        RECT  0.300 164.850 64.700 165.150 ;
        RECT  0.300 165.450 64.700 165.750 ;
        RECT  0.300 166.050 64.700 166.350 ;
        RECT  0.300 166.650 64.700 166.960 ;
        RECT  0.300 167.260 64.700 167.560 ;
        RECT  0.300 167.860 64.700 168.160 ;
        RECT  0.000 169.150 65.000 197.240 ;
        RECT  0.600 0.600 64.400 250.000 ;
        RECT  0.000 198.470 65.000 250.000 ;
        LAYER M2 ;
        RECT  63.180 196.430 63.670 249.400 ;
        RECT  0.600 196.440 64.400 245.485 ;
        RECT  26.530 196.440 64.400 248.790 ;
        RECT  0.600 196.440 22.950 249.400 ;
        RECT  26.530 196.440 27.050 249.400 ;
        RECT  30.390 196.440 64.400 249.400 ;
        RECT  0.600 183.850 64.400 185.680 ;
        RECT  46.230 183.850 51.730 185.870 ;
        RECT  4.895 155.120 7.525 171.290 ;
        RECT  8.170 155.125 8.490 171.290 ;
        RECT  21.080 155.160 21.430 171.290 ;
        RECT  21.730 155.140 22.050 171.290 ;
        RECT  53.655 155.035 53.935 171.290 ;
        RECT  56.365 155.280 56.645 171.290 ;
        RECT  57.120 155.300 57.400 171.290 ;
        RECT  57.835 155.130 58.115 171.290 ;
        RECT  0.600 155.310 64.400 171.290 ;
        RECT  53.895 155.310 55.870 171.370 ;
        RECT  33.190 155.310 33.690 171.375 ;
        RECT  3.210 155.310 3.490 171.380 ;
        RECT  34.655 155.310 38.715 171.480 ;
        RECT  39.605 155.310 42.020 171.480 ;
        RECT  2.000 0.000 63.000 60.210 ;
        RECT  0.600 0.600 64.400 60.210 ;
        RECT  0.600 0.600 1.210 135.520 ;
        RECT  0.600 91.020 64.400 135.520 ;
        RECT  4.080 91.020 60.940 135.690 ;
        RECT  62.580 91.020 62.995 135.710 ;
        LAYER M3 ;
        RECT  0.600 247.660 23.220 248.740 ;
        RECT  0.600 247.660 22.900 249.400 ;
        RECT  26.260 247.660 64.400 248.740 ;
        RECT  26.580 247.660 27.000 249.400 ;
        RECT  30.440 247.660 64.400 249.400 ;
        RECT  0.600 124.090 64.400 129.850 ;
        RECT  1.640 124.090 63.600 135.790 ;
        RECT  1.810 124.090 2.830 154.520 ;
        RECT  3.110 124.090 63.600 171.560 ;
        RECT  4.040 123.970 60.900 171.560 ;
        RECT  1.640 155.040 63.600 171.560 ;
        RECT  1.640 183.580 63.600 185.950 ;
        RECT  5.510 124.090 63.600 200.820 ;
        RECT  1.640 196.170 63.600 200.820 ;
        RECT  0.600 0.600 64.400 60.480 ;
        RECT  2.000 0.000 63.000 88.700 ;
        RECT  0.600 0.600 1.480 91.220 ;
        RECT  0.600 90.750 64.400 91.220 ;
        LAYER TOP_M ;
        RECT  0.600 247.690 64.400 248.850 ;
        RECT  0.600 247.690 23.010 249.400 ;
        RECT  26.470 247.690 27.110 249.400 ;
        RECT  30.330 247.690 64.400 249.400 ;
        RECT  2.000 0.000 63.000 91.190 ;
        RECT  0.600 0.600 64.400 91.190 ;
    END
END pc3t03u

MACRO pc3t03d
    CLASS PAD ;
    FOREIGN pc3t03d 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 65.000 BY 250.000 ;
    SYMMETRY X Y R90 ;
    SITE IOSite_c ;
    PIN PAD
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 55.440  LAYER TOP_M  ;
        ANTENNAPARTIALMETALSIDEAREA 287.938  LAYER M3  ;
        ANTENNAPARTIALMETALSIDEAREA 480.740  LAYER M2  ;
        ANTENNADIFFAREA 2657.280  LAYER TOP_M  ;
        ANTENNADIFFAREA 2657.280  LAYER M3  ;
        ANTENNADIFFAREA 1209.600  LAYER M2  ;
        ANTENNAPARTIALCUTAREA 632.318  LAYER TOP_V  ;
        ANTENNAPARTIALCUTAREA 349.898  LAYER V3  ;
        ANTENNAPARTIALCUTAREA 255.798  LAYER V2  ;
        PORT
        LAYER M3 ;
        RECT  23.740 249.580 25.740 250.000 ;
        LAYER M2 ;
        RECT  2.000 61.000 63.000 90.230 ;
        RECT  23.740 246.275 25.740 250.000 ;
        END
    END PAD
    PIN OEN
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 81.726  LAYER M2  ;
        ANTENNAPARTIALMETALSIDEAREA 67.374  LAYER M1  ;
        ANTENNAPARTIALMETALSIDEAREA 41.679  LAYER M3  ;
        ANTENNADIFFAREA 0.250  LAYER M3  ;
        ANTENNAPARTIALCUTAREA 0.203  LAYER V2  ;
        ANTENNAPARTIALCUTAREA 0.135  LAYER V3  ;
        ANTENNAGATEAREA 8.100  LAYER M2  ;
        ANTENNAGATEAREA 9.900  LAYER M3  ;
        PORT
        LAYER M3 ;
        RECT  28.870 249.580 29.600 250.000 ;
        LAYER M2 ;
        RECT  28.870 249.580 29.600 250.000 ;
        END
    END OEN
    PIN I
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 67.374  LAYER M1  ;
        ANTENNAPARTIALMETALSIDEAREA 80.804  LAYER M2  ;
        ANTENNAPARTIALMETALSIDEAREA 41.096  LAYER M3  ;
        ANTENNADIFFAREA 0.250  LAYER M3  ;
        ANTENNAPARTIALCUTAREA 0.270  LAYER V2  ;
        ANTENNAPARTIALCUTAREA 0.135  LAYER V3  ;
        ANTENNAGATEAREA 18.900  LAYER M2  ;
        ANTENNAGATEAREA 20.700  LAYER M3  ;
        PORT
        LAYER M3 ;
        RECT  27.840 249.580 28.570 250.000 ;
        LAYER M2 ;
        RECT  27.840 249.580 28.570 250.000 ;
        END
    END I
    PIN VDDO
        DIRECTION INOUT ;
        USE power ;
        PORT
        LAYER M3 ;
        RECT  64.200 192.330 65.000 200.640 ;
        RECT  0.000 201.660 65.000 221.520 ;
        RECT  0.000 222.720 65.000 246.820 ;
        RECT  0.000 192.330 0.800 200.640 ;
        LAYER M2 ;
        RECT  0.000 186.470 65.000 195.650 ;
        LAYER TOP_M ;
        RECT  0.000 195.170 65.000 200.640 ;
        RECT  0.000 201.660 65.000 221.520 ;
        RECT  0.000 222.720 65.000 246.820 ;
        END
    END VDDO
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        PORT
        LAYER M3 ;
        RECT  64.200 163.510 65.000 190.890 ;
        RECT  0.000 163.510 0.800 190.890 ;
        LAYER M2 ;
        RECT  0.000 172.080 65.000 183.060 ;
        LAYER TOP_M ;
        RECT  0.000 163.500 65.000 194.560 ;
        END
    END VDD
    PIN VSSO
        DIRECTION INOUT ;
        USE ground ;
        PORT
        LAYER M3 ;
        RECT  0.000 92.060 65.000 123.250 ;
        RECT  64.200 149.940 65.000 162.610 ;
        RECT  0.000 149.940 0.800 162.610 ;
        LAYER M2 ;
        RECT  0.000 147.040 65.000 154.520 ;
        LAYER TOP_M ;
        RECT  0.000 92.060 65.000 123.250 ;
        RECT  0.000 155.410 65.000 162.610 ;
        END
    END VSSO
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        PORT
        LAYER M3 ;
        RECT  64.200 130.690 65.000 148.880 ;
        RECT  0.000 130.690 0.800 148.880 ;
        LAYER M2 ;
        RECT  0.000 136.310 65.000 146.340 ;
        LAYER TOP_M ;
        RECT  0.000 123.850 65.000 154.560 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  2.000 0.000 63.000 250.000 ;
        RECT  0.000 88.990 65.000 130.360 ;
        RECT  0.000 136.510 65.000 157.550 ;
        RECT  0.315 158.150 64.700 158.460 ;
        RECT  0.300 158.930 64.700 159.230 ;
        RECT  0.300 159.530 64.700 159.830 ;
        RECT  0.300 160.130 64.700 160.430 ;
        RECT  0.300 160.730 64.700 161.030 ;
        RECT  0.300 161.330 64.700 161.630 ;
        RECT  0.300 161.910 64.700 162.190 ;
        RECT  0.300 162.490 64.700 162.770 ;
        RECT  0.300 163.070 64.700 163.350 ;
        RECT  0.300 163.650 64.700 163.950 ;
        RECT  0.300 164.250 64.700 164.550 ;
        RECT  0.300 164.850 64.700 165.150 ;
        RECT  0.300 165.450 64.700 165.750 ;
        RECT  0.300 166.050 64.700 166.350 ;
        RECT  0.300 166.650 64.700 166.960 ;
        RECT  0.300 167.260 64.700 167.560 ;
        RECT  0.300 167.860 64.700 168.160 ;
        RECT  0.000 169.150 65.000 197.240 ;
        RECT  0.600 0.600 64.400 250.000 ;
        RECT  0.000 198.470 65.000 250.000 ;
        LAYER M2 ;
        RECT  63.180 196.430 63.670 249.400 ;
        RECT  0.600 196.440 64.400 245.485 ;
        RECT  26.530 196.440 64.400 248.790 ;
        RECT  0.600 196.440 22.950 249.400 ;
        RECT  26.530 196.440 27.050 249.400 ;
        RECT  30.390 196.440 64.400 249.400 ;
        RECT  0.600 183.850 64.400 185.680 ;
        RECT  46.230 183.850 51.730 185.870 ;
        RECT  4.895 155.120 7.525 171.290 ;
        RECT  8.170 155.125 8.490 171.290 ;
        RECT  21.080 155.160 21.430 171.290 ;
        RECT  21.730 155.140 22.050 171.290 ;
        RECT  49.115 155.130 51.355 171.290 ;
        RECT  52.295 155.300 52.605 171.290 ;
        RECT  53.655 155.035 53.935 171.290 ;
        RECT  56.365 155.280 56.645 171.290 ;
        RECT  57.120 155.300 57.400 171.290 ;
        RECT  57.835 155.130 58.115 171.290 ;
        RECT  0.600 155.310 64.400 171.290 ;
        RECT  53.895 155.310 55.870 171.370 ;
        RECT  3.210 155.310 3.490 171.380 ;
        RECT  34.655 155.310 38.715 171.480 ;
        RECT  39.605 155.310 42.020 171.480 ;
        RECT  2.000 0.000 63.000 60.210 ;
        RECT  0.600 0.600 64.400 60.210 ;
        RECT  0.600 0.600 1.210 135.520 ;
        RECT  0.600 91.020 64.400 135.520 ;
        RECT  4.080 91.020 60.940 135.690 ;
        RECT  62.580 91.020 62.995 135.710 ;
        LAYER M3 ;
        RECT  0.600 247.660 23.220 248.740 ;
        RECT  0.600 247.660 22.900 249.400 ;
        RECT  26.260 247.660 64.400 248.740 ;
        RECT  26.580 247.660 27.000 249.400 ;
        RECT  30.440 247.660 64.400 249.400 ;
        RECT  0.600 124.090 64.400 129.850 ;
        RECT  1.640 124.090 63.600 135.790 ;
        RECT  1.810 124.090 2.830 154.520 ;
        RECT  3.110 124.090 63.600 171.560 ;
        RECT  4.040 123.970 60.900 171.560 ;
        RECT  1.640 155.040 63.600 171.560 ;
        RECT  1.640 183.580 63.600 185.950 ;
        RECT  5.510 124.090 63.600 200.820 ;
        RECT  1.640 196.170 63.600 200.820 ;
        RECT  0.600 0.600 64.400 60.480 ;
        RECT  2.000 0.000 63.000 88.700 ;
        RECT  0.600 0.600 1.480 91.220 ;
        RECT  0.600 90.750 64.400 91.220 ;
        LAYER TOP_M ;
        RECT  0.600 247.690 64.400 248.850 ;
        RECT  0.600 247.690 23.010 249.400 ;
        RECT  26.470 247.690 27.110 249.400 ;
        RECT  30.330 247.690 64.400 249.400 ;
        RECT  2.000 0.000 63.000 91.190 ;
        RECT  0.600 0.600 64.400 91.190 ;
    END
END pc3t03d

MACRO pc3t03
    CLASS PAD ;
    FOREIGN pc3t03 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 65.000 BY 250.000 ;
    SYMMETRY X Y R90 ;
    SITE IOSite_c ;
    PIN PAD
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 55.440  LAYER TOP_M  ;
        ANTENNAPARTIALMETALSIDEAREA 287.938  LAYER M3  ;
        ANTENNAPARTIALMETALSIDEAREA 480.740  LAYER M2  ;
        ANTENNADIFFAREA 2657.280  LAYER TOP_M  ;
        ANTENNADIFFAREA 2657.280  LAYER M3  ;
        ANTENNADIFFAREA 1209.600  LAYER M2  ;
        ANTENNAPARTIALCUTAREA 632.318  LAYER TOP_V  ;
        ANTENNAPARTIALCUTAREA 349.898  LAYER V3  ;
        ANTENNAPARTIALCUTAREA 255.798  LAYER V2  ;
        PORT
        LAYER M3 ;
        RECT  23.740 249.580 25.740 250.000 ;
        LAYER M2 ;
        RECT  2.000 61.000 63.000 90.230 ;
        RECT  23.740 246.275 25.740 250.000 ;
        END
    END PAD
    PIN OEN
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 67.374  LAYER M1  ;
        ANTENNAPARTIALMETALSIDEAREA 81.726  LAYER M2  ;
        ANTENNAPARTIALMETALSIDEAREA 41.679  LAYER M3  ;
        ANTENNADIFFAREA 0.250  LAYER M3  ;
        ANTENNAPARTIALCUTAREA 0.203  LAYER V2  ;
        ANTENNAPARTIALCUTAREA 0.135  LAYER V3  ;
        ANTENNAGATEAREA 8.100  LAYER M2  ;
        ANTENNAGATEAREA 9.900  LAYER M3  ;
        PORT
        LAYER M3 ;
        RECT  28.870 249.580 29.600 250.000 ;
        LAYER M2 ;
        RECT  28.870 249.580 29.600 250.000 ;
        END
    END OEN
    PIN I
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 67.374  LAYER M1  ;
        ANTENNAPARTIALMETALSIDEAREA 80.804  LAYER M2  ;
        ANTENNAPARTIALMETALSIDEAREA 41.096  LAYER M3  ;
        ANTENNADIFFAREA 0.250  LAYER M3  ;
        ANTENNAPARTIALCUTAREA 0.270  LAYER V2  ;
        ANTENNAPARTIALCUTAREA 0.135  LAYER V3  ;
        ANTENNAGATEAREA 18.900  LAYER M2  ;
        ANTENNAGATEAREA 20.700  LAYER M3  ;
        PORT
        LAYER M3 ;
        RECT  27.840 249.580 28.570 250.000 ;
        LAYER M2 ;
        RECT  27.840 249.580 28.570 250.000 ;
        END
    END I
    PIN VDDO
        DIRECTION INOUT ;
        USE power ;
        PORT
        LAYER M3 ;
        RECT  64.200 192.330 65.000 200.640 ;
        RECT  0.000 201.660 65.000 221.520 ;
        RECT  0.000 222.720 65.000 246.820 ;
        RECT  0.000 192.330 0.800 200.640 ;
        LAYER M2 ;
        RECT  0.000 186.470 65.000 195.650 ;
        LAYER TOP_M ;
        RECT  0.000 195.170 65.000 200.640 ;
        RECT  0.000 201.660 65.000 221.520 ;
        RECT  0.000 222.720 65.000 246.820 ;
        END
    END VDDO
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        PORT
        LAYER M3 ;
        RECT  64.200 163.510 65.000 190.890 ;
        RECT  0.000 163.510 0.800 190.890 ;
        LAYER M2 ;
        RECT  0.000 172.080 65.000 183.060 ;
        LAYER TOP_M ;
        RECT  0.000 163.500 65.000 194.560 ;
        END
    END VDD
    PIN VSSO
        DIRECTION INOUT ;
        USE ground ;
        PORT
        LAYER M3 ;
        RECT  0.000 92.060 65.000 123.250 ;
        RECT  64.200 149.940 65.000 162.610 ;
        RECT  0.000 149.940 0.800 162.610 ;
        LAYER M2 ;
        RECT  0.000 147.040 65.000 154.520 ;
        LAYER TOP_M ;
        RECT  0.000 92.060 65.000 123.250 ;
        RECT  0.000 155.410 65.000 162.610 ;
        END
    END VSSO
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        PORT
        LAYER M3 ;
        RECT  64.200 130.690 65.000 148.880 ;
        RECT  0.000 130.690 0.800 148.880 ;
        LAYER M2 ;
        RECT  0.000 136.310 65.000 146.340 ;
        LAYER TOP_M ;
        RECT  0.000 123.850 65.000 154.560 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  2.000 0.000 63.000 250.000 ;
        RECT  0.000 88.990 65.000 130.360 ;
        RECT  0.000 136.510 65.000 157.550 ;
        RECT  0.315 158.150 64.700 158.460 ;
        RECT  0.300 158.930 64.700 159.230 ;
        RECT  0.300 159.530 64.700 159.830 ;
        RECT  0.300 160.130 64.700 160.430 ;
        RECT  0.300 160.730 64.700 161.030 ;
        RECT  0.300 161.330 64.700 161.630 ;
        RECT  0.300 161.910 64.700 162.190 ;
        RECT  0.300 162.490 64.700 162.770 ;
        RECT  0.300 163.070 64.700 163.350 ;
        RECT  0.300 163.650 64.700 163.950 ;
        RECT  0.300 164.250 64.700 164.550 ;
        RECT  0.300 164.850 64.700 165.150 ;
        RECT  0.300 165.450 64.700 165.750 ;
        RECT  0.300 166.050 64.700 166.350 ;
        RECT  0.300 166.650 64.700 166.960 ;
        RECT  0.300 167.260 64.700 167.560 ;
        RECT  0.300 167.860 64.700 168.160 ;
        RECT  0.000 169.150 65.000 197.240 ;
        RECT  0.600 0.600 64.400 250.000 ;
        RECT  0.000 198.470 65.000 250.000 ;
        LAYER M2 ;
        RECT  63.180 196.430 63.670 249.400 ;
        RECT  0.600 196.440 64.400 245.485 ;
        RECT  26.530 196.440 64.400 248.790 ;
        RECT  0.600 196.440 22.950 249.400 ;
        RECT  26.530 196.440 27.050 249.400 ;
        RECT  30.390 196.440 64.400 249.400 ;
        RECT  0.600 183.850 64.400 185.680 ;
        RECT  46.230 183.850 51.730 185.870 ;
        RECT  4.895 155.120 7.525 171.290 ;
        RECT  8.170 155.125 8.490 171.290 ;
        RECT  21.080 155.160 21.430 171.290 ;
        RECT  21.730 155.140 22.050 171.290 ;
        RECT  53.655 155.035 53.935 171.290 ;
        RECT  56.365 155.280 56.645 171.290 ;
        RECT  57.120 155.300 57.400 171.290 ;
        RECT  57.835 155.130 58.115 171.290 ;
        RECT  0.600 155.310 64.400 171.290 ;
        RECT  53.895 155.310 55.870 171.370 ;
        RECT  3.210 155.310 3.490 171.380 ;
        RECT  34.655 155.310 38.715 171.480 ;
        RECT  39.605 155.310 42.020 171.480 ;
        RECT  2.000 0.000 63.000 60.210 ;
        RECT  0.600 0.600 64.400 60.210 ;
        RECT  0.600 0.600 1.210 135.520 ;
        RECT  0.600 91.020 64.400 135.520 ;
        RECT  4.080 91.020 60.940 135.690 ;
        RECT  62.580 91.020 62.995 135.710 ;
        LAYER M3 ;
        RECT  0.600 247.660 23.220 248.740 ;
        RECT  0.600 247.660 22.900 249.400 ;
        RECT  26.260 247.660 64.400 248.740 ;
        RECT  26.580 247.660 27.000 249.400 ;
        RECT  30.440 247.660 64.400 249.400 ;
        RECT  0.600 124.090 64.400 129.850 ;
        RECT  1.640 124.090 63.600 135.790 ;
        RECT  1.810 124.090 2.830 154.520 ;
        RECT  3.110 124.090 63.600 171.560 ;
        RECT  4.040 123.970 60.900 171.560 ;
        RECT  1.640 155.040 63.600 171.560 ;
        RECT  1.640 183.580 63.600 185.950 ;
        RECT  5.510 124.090 63.600 200.820 ;
        RECT  1.640 196.170 63.600 200.820 ;
        RECT  0.600 0.600 64.400 60.480 ;
        RECT  2.000 0.000 63.000 88.700 ;
        RECT  0.600 0.600 1.480 91.220 ;
        RECT  0.600 90.750 64.400 91.220 ;
        LAYER TOP_M ;
        RECT  0.600 247.690 64.400 248.850 ;
        RECT  0.600 247.690 23.010 249.400 ;
        RECT  26.470 247.690 27.110 249.400 ;
        RECT  30.330 247.690 64.400 249.400 ;
        RECT  2.000 0.000 63.000 91.190 ;
        RECT  0.600 0.600 64.400 91.190 ;
    END
END pc3t03

MACRO pc3t02u
    CLASS PAD ;
    FOREIGN pc3t02u 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 65.000 BY 250.000 ;
    SYMMETRY X Y R90 ;
    SITE IOSite_c ;
    PIN PAD
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 55.440  LAYER TOP_M  ;
        ANTENNAPARTIALMETALSIDEAREA 287.938  LAYER M3  ;
        ANTENNAPARTIALMETALSIDEAREA 480.740  LAYER M2  ;
        ANTENNADIFFAREA 2657.280  LAYER TOP_M  ;
        ANTENNADIFFAREA 2657.280  LAYER M3  ;
        ANTENNADIFFAREA 1209.600  LAYER M2  ;
        ANTENNAPARTIALCUTAREA 632.318  LAYER TOP_V  ;
        ANTENNAPARTIALCUTAREA 349.898  LAYER V3  ;
        ANTENNAPARTIALCUTAREA 255.798  LAYER V2  ;
        PORT
        LAYER M3 ;
        RECT  23.740 249.580 25.740 250.000 ;
        LAYER M2 ;
        RECT  2.000 61.000 63.000 90.230 ;
        RECT  23.740 246.275 25.740 250.000 ;
        END
    END PAD
    PIN OEN
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 81.726  LAYER M2  ;
        ANTENNAPARTIALMETALSIDEAREA 67.374  LAYER M1  ;
        ANTENNAPARTIALMETALSIDEAREA 41.679  LAYER M3  ;
        ANTENNADIFFAREA 0.250  LAYER M3  ;
        ANTENNAPARTIALCUTAREA 0.203  LAYER V2  ;
        ANTENNAPARTIALCUTAREA 0.135  LAYER V3  ;
        ANTENNAGATEAREA 8.100  LAYER M2  ;
        ANTENNAGATEAREA 9.900  LAYER M3  ;
        PORT
        LAYER M3 ;
        RECT  28.870 249.580 29.600 250.000 ;
        LAYER M2 ;
        RECT  28.870 249.580 29.600 250.000 ;
        END
    END OEN
    PIN I
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 67.374  LAYER M1  ;
        ANTENNAPARTIALMETALSIDEAREA 80.804  LAYER M2  ;
        ANTENNAPARTIALMETALSIDEAREA 41.096  LAYER M3  ;
        ANTENNADIFFAREA 0.250  LAYER M3  ;
        ANTENNAPARTIALCUTAREA 0.270  LAYER V2  ;
        ANTENNAPARTIALCUTAREA 0.135  LAYER V3  ;
        ANTENNAGATEAREA 18.900  LAYER M2  ;
        ANTENNAGATEAREA 20.700  LAYER M3  ;
        PORT
        LAYER M3 ;
        RECT  27.840 249.580 28.570 250.000 ;
        LAYER M2 ;
        RECT  27.840 249.580 28.570 250.000 ;
        END
    END I
    PIN VDDO
        DIRECTION INOUT ;
        USE power ;
        PORT
        LAYER M3 ;
        RECT  64.200 192.330 65.000 200.640 ;
        RECT  0.000 201.660 65.000 221.520 ;
        RECT  0.000 222.720 65.000 246.820 ;
        RECT  0.000 192.330 0.800 200.640 ;
        LAYER M2 ;
        RECT  0.000 186.470 65.000 195.650 ;
        LAYER TOP_M ;
        RECT  0.000 195.170 65.000 200.640 ;
        RECT  0.000 201.660 65.000 221.520 ;
        RECT  0.000 222.720 65.000 246.820 ;
        END
    END VDDO
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        PORT
        LAYER M3 ;
        RECT  64.200 163.510 65.000 190.890 ;
        RECT  0.000 163.510 0.800 190.890 ;
        LAYER M2 ;
        RECT  0.000 172.080 65.000 183.060 ;
        LAYER TOP_M ;
        RECT  0.000 163.500 65.000 194.560 ;
        END
    END VDD
    PIN VSSO
        DIRECTION INOUT ;
        USE ground ;
        PORT
        LAYER M3 ;
        RECT  0.000 92.060 65.000 123.250 ;
        RECT  64.200 149.940 65.000 162.610 ;
        RECT  0.000 149.940 0.800 162.610 ;
        LAYER M2 ;
        RECT  0.000 147.040 65.000 154.520 ;
        LAYER TOP_M ;
        RECT  0.000 92.060 65.000 123.250 ;
        RECT  0.000 155.410 65.000 162.610 ;
        END
    END VSSO
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        PORT
        LAYER M3 ;
        RECT  64.200 130.690 65.000 148.880 ;
        RECT  0.000 130.690 0.800 148.880 ;
        LAYER M2 ;
        RECT  0.000 136.310 65.000 146.340 ;
        LAYER TOP_M ;
        RECT  0.000 123.850 65.000 154.560 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  2.000 0.000 63.000 250.000 ;
        RECT  0.000 88.990 65.000 130.360 ;
        RECT  0.000 136.510 65.000 157.550 ;
        RECT  0.315 158.150 64.700 158.460 ;
        RECT  0.300 158.930 64.700 159.230 ;
        RECT  0.300 159.530 64.700 159.830 ;
        RECT  0.300 160.130 64.700 160.430 ;
        RECT  0.300 160.730 64.700 161.030 ;
        RECT  0.300 161.330 64.700 161.630 ;
        RECT  0.300 161.910 64.700 162.190 ;
        RECT  0.300 162.490 64.700 162.770 ;
        RECT  0.300 163.070 64.700 163.350 ;
        RECT  0.300 163.650 64.700 163.950 ;
        RECT  0.300 164.250 64.700 164.550 ;
        RECT  0.300 164.850 64.700 165.150 ;
        RECT  0.300 165.450 64.700 165.750 ;
        RECT  0.300 166.050 64.700 166.350 ;
        RECT  0.300 166.650 64.700 166.960 ;
        RECT  0.300 167.260 64.700 167.560 ;
        RECT  0.300 167.860 64.700 168.160 ;
        RECT  0.000 169.150 65.000 197.240 ;
        RECT  0.600 0.600 64.400 250.000 ;
        RECT  0.000 198.470 65.000 250.000 ;
        LAYER M2 ;
        RECT  63.180 196.430 63.670 249.400 ;
        RECT  0.600 196.440 64.400 245.485 ;
        RECT  26.530 196.440 64.400 248.790 ;
        RECT  0.600 196.440 22.950 249.400 ;
        RECT  26.530 196.440 27.050 249.400 ;
        RECT  30.390 196.440 64.400 249.400 ;
        RECT  0.600 183.850 64.400 185.680 ;
        RECT  46.230 183.850 51.730 185.870 ;
        RECT  9.050 155.125 9.370 171.290 ;
        RECT  20.490 155.160 20.840 171.290 ;
        RECT  21.140 155.140 21.460 171.290 ;
        RECT  53.655 155.035 53.935 171.290 ;
        RECT  56.365 155.280 56.645 171.290 ;
        RECT  57.120 155.300 57.400 171.290 ;
        RECT  57.835 155.130 58.115 171.290 ;
        RECT  0.600 155.310 64.400 171.290 ;
        RECT  32.465 155.310 32.965 171.370 ;
        RECT  53.895 155.310 55.870 171.370 ;
        RECT  3.225 155.310 3.505 171.380 ;
        RECT  34.655 155.310 38.715 171.480 ;
        RECT  39.605 155.310 42.020 171.480 ;
        RECT  2.000 0.000 63.000 60.210 ;
        RECT  0.600 0.600 64.400 60.210 ;
        RECT  0.600 0.600 1.210 135.520 ;
        RECT  0.600 91.020 64.400 135.520 ;
        RECT  4.080 91.020 60.940 135.690 ;
        RECT  62.580 91.020 62.995 135.710 ;
        LAYER M3 ;
        RECT  0.600 247.660 23.220 248.740 ;
        RECT  0.600 247.660 22.900 249.400 ;
        RECT  26.260 247.660 64.400 248.740 ;
        RECT  26.580 247.660 27.000 249.400 ;
        RECT  30.440 247.660 64.400 249.400 ;
        RECT  0.600 124.090 64.400 129.850 ;
        RECT  1.640 124.090 63.600 135.790 ;
        RECT  1.810 124.090 2.830 154.520 ;
        RECT  3.110 124.090 63.600 171.560 ;
        RECT  4.040 123.970 60.900 171.560 ;
        RECT  1.640 155.040 63.600 171.560 ;
        RECT  1.640 183.580 63.600 185.950 ;
        RECT  5.490 124.090 63.600 200.820 ;
        RECT  1.640 196.170 63.600 200.820 ;
        RECT  0.600 0.600 64.400 60.480 ;
        RECT  2.000 0.000 63.000 88.700 ;
        RECT  0.600 0.600 1.480 91.220 ;
        RECT  0.600 90.750 64.400 91.220 ;
        LAYER TOP_M ;
        RECT  0.600 247.690 64.400 248.850 ;
        RECT  0.600 247.690 23.010 249.400 ;
        RECT  26.470 247.690 27.110 249.400 ;
        RECT  30.330 247.690 64.400 249.400 ;
        RECT  2.000 0.000 63.000 91.190 ;
        RECT  0.600 0.600 64.400 91.190 ;
    END
END pc3t02u

MACRO pc3t02d
    CLASS PAD ;
    FOREIGN pc3t02d 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 65.000 BY 250.000 ;
    SYMMETRY X Y R90 ;
    SITE IOSite_c ;
    PIN PAD
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 55.440  LAYER TOP_M  ;
        ANTENNAPARTIALMETALSIDEAREA 287.938  LAYER M3  ;
        ANTENNAPARTIALMETALSIDEAREA 480.740  LAYER M2  ;
        ANTENNADIFFAREA 2657.280  LAYER TOP_M  ;
        ANTENNADIFFAREA 2657.280  LAYER M3  ;
        ANTENNADIFFAREA 1209.600  LAYER M2  ;
        ANTENNAPARTIALCUTAREA 632.318  LAYER TOP_V  ;
        ANTENNAPARTIALCUTAREA 349.898  LAYER V3  ;
        ANTENNAPARTIALCUTAREA 255.798  LAYER V2  ;
        PORT
        LAYER M3 ;
        RECT  23.740 249.580 25.740 250.000 ;
        LAYER M2 ;
        RECT  2.000 61.000 63.000 90.230 ;
        RECT  23.740 246.275 25.740 250.000 ;
        END
    END PAD
    PIN OEN
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 67.374  LAYER M1  ;
        ANTENNAPARTIALMETALSIDEAREA 81.726  LAYER M2  ;
        ANTENNAPARTIALMETALSIDEAREA 41.679  LAYER M3  ;
        ANTENNADIFFAREA 0.250  LAYER M3  ;
        ANTENNAPARTIALCUTAREA 0.203  LAYER V2  ;
        ANTENNAPARTIALCUTAREA 0.135  LAYER V3  ;
        ANTENNAGATEAREA 8.100  LAYER M2  ;
        ANTENNAGATEAREA 9.900  LAYER M3  ;
        PORT
        LAYER M3 ;
        RECT  28.870 249.580 29.600 250.000 ;
        LAYER M2 ;
        RECT  28.870 249.580 29.600 250.000 ;
        END
    END OEN
    PIN I
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 80.804  LAYER M2  ;
        ANTENNAPARTIALMETALSIDEAREA 67.374  LAYER M1  ;
        ANTENNAPARTIALMETALSIDEAREA 41.096  LAYER M3  ;
        ANTENNADIFFAREA 0.250  LAYER M3  ;
        ANTENNAPARTIALCUTAREA 0.135  LAYER V3  ;
        ANTENNAPARTIALCUTAREA 0.270  LAYER V2  ;
        ANTENNAGATEAREA 18.900  LAYER M2  ;
        ANTENNAGATEAREA 20.700  LAYER M3  ;
        PORT
        LAYER M3 ;
        RECT  27.840 249.580 28.570 250.000 ;
        LAYER M2 ;
        RECT  27.840 249.580 28.570 250.000 ;
        END
    END I
    PIN VDDO
        DIRECTION INOUT ;
        USE power ;
        PORT
        LAYER M3 ;
        RECT  64.200 192.330 65.000 200.640 ;
        RECT  0.000 201.660 65.000 221.520 ;
        RECT  0.000 222.720 65.000 246.820 ;
        RECT  0.000 192.330 0.800 200.640 ;
        LAYER M2 ;
        RECT  0.000 186.470 65.000 195.650 ;
        LAYER TOP_M ;
        RECT  0.000 195.170 65.000 200.640 ;
        RECT  0.000 201.660 65.000 221.520 ;
        RECT  0.000 222.720 65.000 246.820 ;
        END
    END VDDO
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        PORT
        LAYER M3 ;
        RECT  64.200 163.510 65.000 190.890 ;
        RECT  0.000 163.510 0.800 190.890 ;
        LAYER M2 ;
        RECT  0.000 172.080 65.000 183.060 ;
        LAYER TOP_M ;
        RECT  0.000 163.500 65.000 194.560 ;
        END
    END VDD
    PIN VSSO
        DIRECTION INOUT ;
        USE ground ;
        PORT
        LAYER M3 ;
        RECT  0.000 92.060 65.000 123.250 ;
        RECT  64.200 149.940 65.000 162.610 ;
        RECT  0.000 149.940 0.800 162.610 ;
        LAYER M2 ;
        RECT  0.000 147.040 65.000 154.520 ;
        LAYER TOP_M ;
        RECT  0.000 92.060 65.000 123.250 ;
        RECT  0.000 155.410 65.000 162.610 ;
        END
    END VSSO
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        PORT
        LAYER M3 ;
        RECT  64.200 130.690 65.000 148.880 ;
        RECT  0.000 130.690 0.800 148.880 ;
        LAYER M2 ;
        RECT  0.000 136.310 65.000 146.340 ;
        LAYER TOP_M ;
        RECT  0.000 123.850 65.000 154.560 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  2.000 0.000 63.000 250.000 ;
        RECT  0.000 88.990 65.000 130.360 ;
        RECT  0.000 136.510 65.000 157.550 ;
        RECT  0.315 158.150 64.700 158.460 ;
        RECT  0.300 158.930 64.700 159.230 ;
        RECT  0.300 159.530 64.700 159.830 ;
        RECT  0.300 160.130 64.700 160.430 ;
        RECT  0.300 160.730 64.700 161.030 ;
        RECT  0.300 161.330 64.700 161.630 ;
        RECT  0.300 161.910 64.700 162.190 ;
        RECT  0.300 162.490 64.700 162.770 ;
        RECT  0.300 163.070 64.700 163.350 ;
        RECT  0.300 163.650 64.700 163.950 ;
        RECT  0.300 164.250 64.700 164.550 ;
        RECT  0.300 164.850 64.700 165.150 ;
        RECT  0.300 165.450 64.700 165.750 ;
        RECT  0.300 166.050 64.700 166.350 ;
        RECT  0.300 166.650 64.700 166.960 ;
        RECT  0.300 167.260 64.700 167.560 ;
        RECT  0.300 167.860 64.700 168.160 ;
        RECT  0.000 169.150 65.000 197.240 ;
        RECT  0.600 0.600 64.400 250.000 ;
        RECT  0.000 198.470 65.000 250.000 ;
        LAYER M2 ;
        RECT  63.180 196.430 63.670 249.400 ;
        RECT  0.600 196.440 64.400 245.485 ;
        RECT  26.530 196.440 64.400 248.790 ;
        RECT  0.600 196.440 22.950 249.400 ;
        RECT  26.530 196.440 27.050 249.400 ;
        RECT  30.390 196.440 64.400 249.400 ;
        RECT  0.600 183.850 64.400 185.680 ;
        RECT  46.230 183.850 51.730 185.870 ;
        RECT  9.050 155.125 9.370 171.290 ;
        RECT  20.490 155.160 20.840 171.290 ;
        RECT  21.140 155.140 21.460 171.290 ;
        RECT  49.270 155.135 51.510 171.290 ;
        RECT  52.450 155.305 52.760 171.290 ;
        RECT  53.655 155.035 53.935 171.290 ;
        RECT  56.365 155.280 56.645 171.290 ;
        RECT  57.120 155.300 57.400 171.290 ;
        RECT  57.835 155.130 58.115 171.290 ;
        RECT  0.600 155.310 64.400 171.290 ;
        RECT  53.895 155.310 55.870 171.370 ;
        RECT  3.225 155.310 3.505 171.380 ;
        RECT  34.655 155.310 38.715 171.480 ;
        RECT  39.605 155.310 42.020 171.480 ;
        RECT  2.000 0.000 63.000 60.210 ;
        RECT  0.600 0.600 64.400 60.210 ;
        RECT  0.600 0.600 1.210 135.520 ;
        RECT  0.600 91.020 64.400 135.520 ;
        RECT  4.080 91.020 60.940 135.690 ;
        RECT  62.580 91.020 62.995 135.710 ;
        LAYER M3 ;
        RECT  0.600 247.660 23.220 248.740 ;
        RECT  0.600 247.660 22.900 249.400 ;
        RECT  26.260 247.660 64.400 248.740 ;
        RECT  26.580 247.660 27.000 249.400 ;
        RECT  30.440 247.660 64.400 249.400 ;
        RECT  0.600 124.090 64.400 129.850 ;
        RECT  1.640 124.090 63.600 135.790 ;
        RECT  1.810 124.090 2.830 154.520 ;
        RECT  3.110 124.090 63.600 171.560 ;
        RECT  4.040 123.970 60.900 171.560 ;
        RECT  1.640 155.040 63.600 171.560 ;
        RECT  1.640 183.580 63.600 185.950 ;
        RECT  5.490 124.090 63.600 200.820 ;
        RECT  1.640 196.170 63.600 200.820 ;
        RECT  0.600 0.600 64.400 60.480 ;
        RECT  2.000 0.000 63.000 88.700 ;
        RECT  0.600 0.600 1.480 91.220 ;
        RECT  0.600 90.750 64.400 91.220 ;
        LAYER TOP_M ;
        RECT  0.600 247.690 64.400 248.850 ;
        RECT  0.600 247.690 23.010 249.400 ;
        RECT  26.470 247.690 27.110 249.400 ;
        RECT  30.330 247.690 64.400 249.400 ;
        RECT  2.000 0.000 63.000 91.190 ;
        RECT  0.600 0.600 64.400 91.190 ;
    END
END pc3t02d

MACRO pc3t02
    CLASS PAD ;
    FOREIGN pc3t02 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 65.000 BY 250.000 ;
    SYMMETRY X Y R90 ;
    SITE IOSite_c ;
    PIN PAD
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 55.440  LAYER TOP_M  ;
        ANTENNAPARTIALMETALSIDEAREA 287.938  LAYER M3  ;
        ANTENNAPARTIALMETALSIDEAREA 480.740  LAYER M2  ;
        ANTENNADIFFAREA 2657.280  LAYER TOP_M  ;
        ANTENNADIFFAREA 2657.280  LAYER M3  ;
        ANTENNADIFFAREA 1209.600  LAYER M2  ;
        ANTENNAPARTIALCUTAREA 632.318  LAYER TOP_V  ;
        ANTENNAPARTIALCUTAREA 349.898  LAYER V3  ;
        ANTENNAPARTIALCUTAREA 255.798  LAYER V2  ;
        PORT
        LAYER M3 ;
        RECT  23.740 249.580 25.740 250.000 ;
        LAYER M2 ;
        RECT  2.000 61.000 63.000 90.230 ;
        RECT  23.740 246.275 25.740 250.000 ;
        END
    END PAD
    PIN OEN
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 67.374  LAYER M1  ;
        ANTENNAPARTIALMETALSIDEAREA 81.726  LAYER M2  ;
        ANTENNAPARTIALMETALSIDEAREA 41.679  LAYER M3  ;
        ANTENNADIFFAREA 0.250  LAYER M3  ;
        ANTENNAPARTIALCUTAREA 0.203  LAYER V2  ;
        ANTENNAPARTIALCUTAREA 0.135  LAYER V3  ;
        ANTENNAGATEAREA 8.100  LAYER M2  ;
        ANTENNAGATEAREA 9.900  LAYER M3  ;
        PORT
        LAYER M3 ;
        RECT  28.870 249.580 29.600 250.000 ;
        LAYER M2 ;
        RECT  28.870 249.580 29.600 250.000 ;
        END
    END OEN
    PIN I
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 67.374  LAYER M1  ;
        ANTENNAPARTIALMETALSIDEAREA 80.804  LAYER M2  ;
        ANTENNAPARTIALMETALSIDEAREA 41.096  LAYER M3  ;
        ANTENNADIFFAREA 0.250  LAYER M3  ;
        ANTENNAPARTIALCUTAREA 0.270  LAYER V2  ;
        ANTENNAPARTIALCUTAREA 0.135  LAYER V3  ;
        ANTENNAGATEAREA 18.900  LAYER M2  ;
        ANTENNAGATEAREA 20.700  LAYER M3  ;
        PORT
        LAYER M3 ;
        RECT  27.840 249.580 28.570 250.000 ;
        LAYER M2 ;
        RECT  27.840 249.580 28.570 250.000 ;
        END
    END I
    PIN VDDO
        DIRECTION INOUT ;
        USE power ;
        PORT
        LAYER M3 ;
        RECT  64.200 192.330 65.000 200.640 ;
        RECT  0.000 201.660 65.000 221.520 ;
        RECT  0.000 222.720 65.000 246.820 ;
        RECT  0.000 192.330 0.800 200.640 ;
        LAYER M2 ;
        RECT  0.000 186.470 65.000 195.650 ;
        LAYER TOP_M ;
        RECT  0.000 195.170 65.000 200.640 ;
        RECT  0.000 201.660 65.000 221.520 ;
        RECT  0.000 222.720 65.000 246.820 ;
        END
    END VDDO
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        PORT
        LAYER M3 ;
        RECT  64.200 163.510 65.000 190.890 ;
        RECT  0.000 163.510 0.800 190.890 ;
        LAYER M2 ;
        RECT  0.000 172.080 65.000 183.060 ;
        LAYER TOP_M ;
        RECT  0.000 163.500 65.000 194.560 ;
        END
    END VDD
    PIN VSSO
        DIRECTION INOUT ;
        USE ground ;
        PORT
        LAYER M3 ;
        RECT  0.000 92.060 65.000 123.250 ;
        RECT  64.200 149.940 65.000 162.610 ;
        RECT  0.000 149.940 0.800 162.610 ;
        LAYER M2 ;
        RECT  0.000 147.040 65.000 154.520 ;
        LAYER TOP_M ;
        RECT  0.000 92.060 65.000 123.250 ;
        RECT  0.000 155.410 65.000 162.610 ;
        END
    END VSSO
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        PORT
        LAYER M3 ;
        RECT  64.200 130.690 65.000 148.880 ;
        RECT  0.000 130.690 0.800 148.880 ;
        LAYER M2 ;
        RECT  0.000 136.310 65.000 146.340 ;
        LAYER TOP_M ;
        RECT  0.000 123.850 65.000 154.560 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  2.000 0.000 63.000 250.000 ;
        RECT  0.000 88.990 65.000 130.360 ;
        RECT  0.000 136.510 65.000 157.550 ;
        RECT  0.315 158.150 64.700 158.460 ;
        RECT  0.300 158.930 64.700 159.230 ;
        RECT  0.300 159.530 64.700 159.830 ;
        RECT  0.300 160.130 64.700 160.430 ;
        RECT  0.300 160.730 64.700 161.030 ;
        RECT  0.300 161.330 64.700 161.630 ;
        RECT  0.300 161.910 64.700 162.190 ;
        RECT  0.300 162.490 64.700 162.770 ;
        RECT  0.300 163.070 64.700 163.350 ;
        RECT  0.300 163.650 64.700 163.950 ;
        RECT  0.300 164.250 64.700 164.550 ;
        RECT  0.300 164.850 64.700 165.150 ;
        RECT  0.300 165.450 64.700 165.750 ;
        RECT  0.300 166.050 64.700 166.350 ;
        RECT  0.300 166.650 64.700 166.960 ;
        RECT  0.300 167.260 64.700 167.560 ;
        RECT  0.300 167.860 64.700 168.160 ;
        RECT  0.000 169.150 65.000 197.240 ;
        RECT  0.600 0.600 64.400 250.000 ;
        RECT  0.000 198.470 65.000 250.000 ;
        LAYER M2 ;
        RECT  63.180 196.430 63.670 249.400 ;
        RECT  0.600 196.440 64.400 245.485 ;
        RECT  26.530 196.440 64.400 248.790 ;
        RECT  0.600 196.440 22.950 249.400 ;
        RECT  26.530 196.440 27.050 249.400 ;
        RECT  30.390 196.440 64.400 249.400 ;
        RECT  0.600 183.850 64.400 185.680 ;
        RECT  46.230 183.850 51.730 185.870 ;
        RECT  9.050 155.125 9.370 171.290 ;
        RECT  20.490 155.160 20.840 171.290 ;
        RECT  21.140 155.140 21.460 171.290 ;
        RECT  53.655 155.035 53.935 171.290 ;
        RECT  56.365 155.280 56.645 171.290 ;
        RECT  57.120 155.300 57.400 171.290 ;
        RECT  57.835 155.130 58.115 171.290 ;
        RECT  0.600 155.310 64.400 171.290 ;
        RECT  53.895 155.310 55.870 171.370 ;
        RECT  3.225 155.310 3.505 171.380 ;
        RECT  34.655 155.310 38.715 171.480 ;
        RECT  39.605 155.310 42.020 171.480 ;
        RECT  2.000 0.000 63.000 60.210 ;
        RECT  0.600 0.600 64.400 60.210 ;
        RECT  0.600 0.600 1.210 135.520 ;
        RECT  0.600 91.020 64.400 135.520 ;
        RECT  4.080 91.020 60.940 135.690 ;
        RECT  62.580 91.020 62.995 135.710 ;
        LAYER M3 ;
        RECT  0.600 247.660 23.220 248.740 ;
        RECT  0.600 247.660 22.900 249.400 ;
        RECT  26.260 247.660 64.400 248.740 ;
        RECT  26.580 247.660 27.000 249.400 ;
        RECT  30.440 247.660 64.400 249.400 ;
        RECT  0.600 124.090 64.400 129.850 ;
        RECT  1.640 124.090 63.600 135.790 ;
        RECT  1.810 124.090 2.830 154.520 ;
        RECT  3.110 124.090 63.600 171.560 ;
        RECT  4.040 123.970 60.900 171.560 ;
        RECT  1.640 155.040 63.600 171.560 ;
        RECT  1.640 183.580 63.600 185.950 ;
        RECT  5.490 124.090 63.600 200.820 ;
        RECT  1.640 196.170 63.600 200.820 ;
        RECT  0.600 0.600 64.400 60.480 ;
        RECT  2.000 0.000 63.000 88.700 ;
        RECT  0.600 0.600 1.480 91.220 ;
        RECT  0.600 90.750 64.400 91.220 ;
        LAYER TOP_M ;
        RECT  0.600 247.690 64.400 248.850 ;
        RECT  0.600 247.690 23.010 249.400 ;
        RECT  26.470 247.690 27.110 249.400 ;
        RECT  30.330 247.690 64.400 249.400 ;
        RECT  2.000 0.000 63.000 91.190 ;
        RECT  0.600 0.600 64.400 91.190 ;
    END
END pc3t02

MACRO pc3t01u
    CLASS PAD ;
    FOREIGN pc3t01u 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 65.000 BY 250.000 ;
    SYMMETRY X Y R90 ;
    SITE IOSite_c ;
    PIN PAD
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 55.440  LAYER TOP_M  ;
        ANTENNAPARTIALMETALSIDEAREA 287.938  LAYER M3  ;
        ANTENNAPARTIALMETALSIDEAREA 480.740  LAYER M2  ;
        ANTENNADIFFAREA 2657.280  LAYER TOP_M  ;
        ANTENNADIFFAREA 2657.280  LAYER M3  ;
        ANTENNADIFFAREA 1209.600  LAYER M2  ;
        ANTENNAPARTIALCUTAREA 632.318  LAYER TOP_V  ;
        ANTENNAPARTIALCUTAREA 349.898  LAYER V3  ;
        ANTENNAPARTIALCUTAREA 255.798  LAYER V2  ;
        PORT
        LAYER M3 ;
        RECT  23.740 249.580 25.740 250.000 ;
        LAYER M2 ;
        RECT  2.000 61.000 63.000 90.230 ;
        RECT  23.740 246.275 25.740 250.000 ;
        END
    END PAD
    PIN OEN
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 81.726  LAYER M2  ;
        ANTENNAPARTIALMETALSIDEAREA 67.374  LAYER M1  ;
        ANTENNAPARTIALMETALSIDEAREA 41.679  LAYER M3  ;
        ANTENNADIFFAREA 0.250  LAYER M3  ;
        ANTENNAPARTIALCUTAREA 0.203  LAYER V2  ;
        ANTENNAPARTIALCUTAREA 0.135  LAYER V3  ;
        ANTENNAGATEAREA 8.100  LAYER M2  ;
        ANTENNAGATEAREA 9.900  LAYER M3  ;
        PORT
        LAYER M3 ;
        RECT  28.870 249.580 29.600 250.000 ;
        LAYER M2 ;
        RECT  28.870 249.580 29.600 250.000 ;
        END
    END OEN
    PIN I
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 67.374  LAYER M1  ;
        ANTENNAPARTIALMETALSIDEAREA 80.804  LAYER M2  ;
        ANTENNAPARTIALMETALSIDEAREA 41.096  LAYER M3  ;
        ANTENNADIFFAREA 0.250  LAYER M3  ;
        ANTENNAPARTIALCUTAREA 0.203  LAYER V2  ;
        ANTENNAPARTIALCUTAREA 0.135  LAYER V3  ;
        ANTENNAGATEAREA 8.100  LAYER M2  ;
        ANTENNAGATEAREA 9.900  LAYER M3  ;
        PORT
        LAYER M3 ;
        RECT  27.840 249.580 28.570 250.000 ;
        LAYER M2 ;
        RECT  27.840 249.580 28.570 250.000 ;
        END
    END I
    PIN VDDO
        DIRECTION INOUT ;
        USE power ;
        PORT
        LAYER M3 ;
        RECT  64.200 192.330 65.000 200.640 ;
        RECT  0.000 201.660 65.000 221.520 ;
        RECT  0.000 222.720 65.000 246.820 ;
        RECT  0.000 192.330 0.800 200.640 ;
        LAYER M2 ;
        RECT  0.000 186.470 65.000 195.650 ;
        LAYER TOP_M ;
        RECT  0.000 195.170 65.000 200.640 ;
        RECT  0.000 201.660 65.000 221.520 ;
        RECT  0.000 222.720 65.000 246.820 ;
        END
    END VDDO
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        PORT
        LAYER M3 ;
        RECT  64.200 163.510 65.000 190.890 ;
        RECT  0.000 163.510 0.800 190.890 ;
        LAYER M2 ;
        RECT  0.000 172.080 65.000 183.060 ;
        LAYER TOP_M ;
        RECT  0.000 163.500 65.000 194.560 ;
        END
    END VDD
    PIN VSSO
        DIRECTION INOUT ;
        USE ground ;
        PORT
        LAYER M3 ;
        RECT  0.000 92.060 65.000 123.250 ;
        RECT  64.200 149.940 65.000 162.610 ;
        RECT  0.000 149.940 0.800 162.610 ;
        LAYER M2 ;
        RECT  0.000 147.040 65.000 154.520 ;
        LAYER TOP_M ;
        RECT  0.000 92.060 65.000 123.250 ;
        RECT  0.000 155.410 65.000 162.610 ;
        END
    END VSSO
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        PORT
        LAYER M3 ;
        RECT  64.200 130.690 65.000 148.880 ;
        RECT  0.000 130.690 0.800 148.880 ;
        LAYER M2 ;
        RECT  0.000 136.310 65.000 146.340 ;
        LAYER TOP_M ;
        RECT  0.000 123.850 65.000 154.560 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  2.000 0.000 63.000 250.000 ;
        RECT  0.000 88.990 65.000 130.360 ;
        RECT  0.000 136.510 65.000 157.550 ;
        RECT  0.315 158.150 64.700 158.460 ;
        RECT  0.300 158.930 64.700 159.230 ;
        RECT  0.300 159.530 64.700 159.830 ;
        RECT  0.300 160.130 64.700 160.430 ;
        RECT  0.300 160.730 64.700 161.030 ;
        RECT  0.300 161.330 64.700 161.630 ;
        RECT  0.300 161.910 64.700 162.190 ;
        RECT  0.300 162.490 64.700 162.770 ;
        RECT  0.300 163.070 64.700 163.350 ;
        RECT  0.300 163.650 64.700 163.950 ;
        RECT  0.300 164.250 64.700 164.550 ;
        RECT  0.300 164.850 64.700 165.150 ;
        RECT  0.300 165.450 64.700 165.750 ;
        RECT  0.300 166.050 64.700 166.350 ;
        RECT  0.300 166.650 64.700 166.960 ;
        RECT  0.300 167.260 64.700 167.560 ;
        RECT  0.300 167.860 64.700 168.160 ;
        RECT  0.000 169.150 65.000 197.240 ;
        RECT  0.600 0.600 64.400 250.000 ;
        RECT  0.000 198.470 65.000 250.000 ;
        LAYER M2 ;
        RECT  63.180 196.430 63.670 249.400 ;
        RECT  0.600 196.440 64.400 245.485 ;
        RECT  26.530 196.440 64.400 248.790 ;
        RECT  0.600 196.440 22.950 249.400 ;
        RECT  26.530 196.440 27.050 249.400 ;
        RECT  30.390 196.440 64.400 249.400 ;
        RECT  0.600 183.850 64.400 185.680 ;
        RECT  46.230 183.850 51.730 185.870 ;
        RECT  19.790 155.160 20.140 171.290 ;
        RECT  20.440 155.140 20.760 171.290 ;
        RECT  53.655 155.035 53.935 171.290 ;
        RECT  56.365 155.280 56.645 171.290 ;
        RECT  57.120 155.300 57.400 171.290 ;
        RECT  57.835 155.130 58.115 171.290 ;
        RECT  0.600 155.310 64.400 171.290 ;
        RECT  53.895 155.310 55.870 171.370 ;
        RECT  31.780 155.310 32.280 171.375 ;
        RECT  3.210 155.310 3.490 171.380 ;
        RECT  34.655 155.310 38.715 171.480 ;
        RECT  39.605 155.310 42.020 171.480 ;
        RECT  2.000 0.000 63.000 60.210 ;
        RECT  0.600 0.600 64.400 60.210 ;
        RECT  0.600 0.600 1.210 135.520 ;
        RECT  0.600 91.020 64.400 135.520 ;
        RECT  4.080 91.020 60.940 135.690 ;
        RECT  62.580 91.020 62.995 135.710 ;
        LAYER M3 ;
        RECT  0.600 247.660 23.220 248.740 ;
        RECT  0.600 247.660 22.900 249.400 ;
        RECT  26.260 247.660 64.400 248.740 ;
        RECT  26.580 247.660 27.000 249.400 ;
        RECT  30.440 247.660 64.400 249.400 ;
        RECT  0.600 124.090 64.400 129.850 ;
        RECT  3.990 123.970 60.900 135.790 ;
        RECT  1.640 124.090 63.600 135.790 ;
        RECT  1.810 124.090 2.830 154.520 ;
        RECT  5.155 123.970 60.900 171.560 ;
        RECT  1.640 155.040 63.600 171.560 ;
        RECT  1.640 183.580 63.600 185.950 ;
        RECT  5.490 124.090 63.600 200.820 ;
        RECT  1.640 196.170 63.600 200.820 ;
        RECT  0.600 0.600 64.400 60.480 ;
        RECT  2.000 0.000 63.000 88.700 ;
        RECT  0.600 0.600 1.480 91.220 ;
        RECT  0.600 90.750 64.400 91.220 ;
        LAYER TOP_M ;
        RECT  0.600 247.690 64.400 248.850 ;
        RECT  0.600 247.690 23.010 249.400 ;
        RECT  26.470 247.690 27.110 249.400 ;
        RECT  30.330 247.690 64.400 249.400 ;
        RECT  2.000 0.000 63.000 91.190 ;
        RECT  0.600 0.600 64.400 91.190 ;
    END
END pc3t01u

MACRO pc3t01d
    CLASS PAD ;
    FOREIGN pc3t01d 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 65.000 BY 250.000 ;
    SYMMETRY X Y R90 ;
    SITE IOSite_c ;
    PIN PAD
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 55.440  LAYER TOP_M  ;
        ANTENNAPARTIALMETALSIDEAREA 287.938  LAYER M3  ;
        ANTENNAPARTIALMETALSIDEAREA 480.740  LAYER M2  ;
        ANTENNADIFFAREA 2657.280  LAYER TOP_M  ;
        ANTENNADIFFAREA 2657.280  LAYER M3  ;
        ANTENNADIFFAREA 1209.600  LAYER M2  ;
        ANTENNAPARTIALCUTAREA 632.318  LAYER TOP_V  ;
        ANTENNAPARTIALCUTAREA 349.898  LAYER V3  ;
        ANTENNAPARTIALCUTAREA 255.798  LAYER V2  ;
        PORT
        LAYER M3 ;
        RECT  23.740 249.580 25.740 250.000 ;
        LAYER M2 ;
        RECT  2.000 61.000 63.000 90.230 ;
        RECT  23.740 246.275 25.740 250.000 ;
        END
    END PAD
    PIN OEN
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 81.726  LAYER M2  ;
        ANTENNAPARTIALMETALSIDEAREA 67.374  LAYER M1  ;
        ANTENNAPARTIALMETALSIDEAREA 41.679  LAYER M3  ;
        ANTENNADIFFAREA 0.250  LAYER M3  ;
        ANTENNAPARTIALCUTAREA 0.203  LAYER V2  ;
        ANTENNAPARTIALCUTAREA 0.135  LAYER V3  ;
        ANTENNAGATEAREA 8.100  LAYER M2  ;
        ANTENNAGATEAREA 9.900  LAYER M3  ;
        PORT
        LAYER M3 ;
        RECT  28.870 249.580 29.600 250.000 ;
        LAYER M2 ;
        RECT  28.870 249.580 29.600 250.000 ;
        END
    END OEN
    PIN I
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 67.374  LAYER M1  ;
        ANTENNAPARTIALMETALSIDEAREA 80.804  LAYER M2  ;
        ANTENNAPARTIALMETALSIDEAREA 41.096  LAYER M3  ;
        ANTENNADIFFAREA 0.250  LAYER M3  ;
        ANTENNAPARTIALCUTAREA 0.203  LAYER V2  ;
        ANTENNAPARTIALCUTAREA 0.135  LAYER V3  ;
        ANTENNAGATEAREA 8.100  LAYER M2  ;
        ANTENNAGATEAREA 9.900  LAYER M3  ;
        PORT
        LAYER M3 ;
        RECT  27.840 249.580 28.570 250.000 ;
        LAYER M2 ;
        RECT  27.840 249.580 28.570 250.000 ;
        END
    END I
    PIN VDDO
        DIRECTION INOUT ;
        USE power ;
        PORT
        LAYER M3 ;
        RECT  64.200 192.330 65.000 200.640 ;
        RECT  0.000 201.660 65.000 221.520 ;
        RECT  0.000 222.720 65.000 246.820 ;
        RECT  0.000 192.330 0.800 200.640 ;
        LAYER M2 ;
        RECT  0.000 186.470 65.000 195.650 ;
        LAYER TOP_M ;
        RECT  0.000 195.170 65.000 200.640 ;
        RECT  0.000 201.660 65.000 221.520 ;
        RECT  0.000 222.720 65.000 246.820 ;
        END
    END VDDO
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        PORT
        LAYER M3 ;
        RECT  64.200 163.510 65.000 190.890 ;
        RECT  0.000 163.510 0.800 190.890 ;
        LAYER M2 ;
        RECT  0.000 172.080 65.000 183.060 ;
        LAYER TOP_M ;
        RECT  0.000 163.500 65.000 194.560 ;
        END
    END VDD
    PIN VSSO
        DIRECTION INOUT ;
        USE ground ;
        PORT
        LAYER M3 ;
        RECT  0.000 92.060 65.000 123.250 ;
        RECT  64.200 149.940 65.000 162.610 ;
        RECT  0.000 149.940 0.800 162.610 ;
        LAYER M2 ;
        RECT  0.000 147.040 65.000 154.520 ;
        LAYER TOP_M ;
        RECT  0.000 92.060 65.000 123.250 ;
        RECT  0.000 155.410 65.000 162.610 ;
        END
    END VSSO
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        PORT
        LAYER M3 ;
        RECT  64.200 130.690 65.000 148.880 ;
        RECT  0.000 130.690 0.800 148.880 ;
        LAYER M2 ;
        RECT  0.000 136.310 65.000 146.340 ;
        LAYER TOP_M ;
        RECT  0.000 123.850 65.000 154.560 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  2.000 0.000 63.000 250.000 ;
        RECT  0.000 88.990 65.000 130.360 ;
        RECT  0.000 136.510 65.000 157.550 ;
        RECT  0.315 158.150 64.700 158.460 ;
        RECT  0.300 158.930 64.700 159.230 ;
        RECT  0.300 159.530 64.700 159.830 ;
        RECT  0.300 160.130 64.700 160.430 ;
        RECT  0.300 160.730 64.700 161.030 ;
        RECT  0.300 161.330 64.700 161.630 ;
        RECT  0.300 161.910 64.700 162.190 ;
        RECT  0.300 162.490 64.700 162.770 ;
        RECT  0.300 163.070 64.700 163.350 ;
        RECT  0.300 163.650 64.700 163.950 ;
        RECT  0.300 164.250 64.700 164.550 ;
        RECT  0.300 164.850 64.700 165.150 ;
        RECT  0.300 165.450 64.700 165.750 ;
        RECT  0.300 166.050 64.700 166.350 ;
        RECT  0.300 166.650 64.700 166.960 ;
        RECT  0.300 167.260 64.700 167.560 ;
        RECT  0.300 167.860 64.700 168.160 ;
        RECT  0.000 169.150 65.000 197.240 ;
        RECT  0.600 0.600 64.400 250.000 ;
        RECT  0.000 198.470 65.000 250.000 ;
        LAYER M2 ;
        RECT  63.180 196.430 63.670 249.400 ;
        RECT  0.600 196.440 64.400 245.485 ;
        RECT  26.530 196.440 64.400 248.790 ;
        RECT  0.600 196.440 22.950 249.400 ;
        RECT  26.530 196.440 27.050 249.400 ;
        RECT  30.390 196.440 64.400 249.400 ;
        RECT  0.600 183.850 64.400 185.680 ;
        RECT  46.230 183.850 51.730 185.870 ;
        RECT  19.790 155.160 20.140 171.290 ;
        RECT  20.440 155.140 20.760 171.290 ;
        RECT  49.330 155.130 51.570 171.290 ;
        RECT  52.510 155.300 52.820 171.290 ;
        RECT  53.655 155.035 53.935 171.290 ;
        RECT  56.365 155.280 56.645 171.290 ;
        RECT  57.120 155.300 57.400 171.290 ;
        RECT  57.835 155.130 58.115 171.290 ;
        RECT  0.600 155.310 64.400 171.290 ;
        RECT  53.895 155.310 55.870 171.370 ;
        RECT  3.210 155.310 3.490 171.380 ;
        RECT  34.655 155.310 38.715 171.480 ;
        RECT  39.605 155.310 42.020 171.480 ;
        RECT  2.000 0.000 63.000 60.210 ;
        RECT  0.600 0.600 64.400 60.210 ;
        RECT  0.600 0.600 1.210 135.520 ;
        RECT  0.600 91.020 64.400 135.520 ;
        RECT  4.080 91.020 60.940 135.690 ;
        RECT  62.580 91.020 62.995 135.710 ;
        LAYER M3 ;
        RECT  0.600 247.660 23.220 248.740 ;
        RECT  0.600 247.660 22.900 249.400 ;
        RECT  26.260 247.660 64.400 248.740 ;
        RECT  26.580 247.660 27.000 249.400 ;
        RECT  30.440 247.660 64.400 249.400 ;
        RECT  0.600 124.090 64.400 129.850 ;
        RECT  3.990 123.970 60.900 135.790 ;
        RECT  1.640 124.090 63.600 135.790 ;
        RECT  1.810 124.090 2.830 154.520 ;
        RECT  5.155 123.970 60.900 171.560 ;
        RECT  1.640 155.040 63.600 171.560 ;
        RECT  1.640 183.580 63.600 185.950 ;
        RECT  5.490 124.090 63.600 200.820 ;
        RECT  1.640 196.170 63.600 200.820 ;
        RECT  0.600 0.600 64.400 60.480 ;
        RECT  2.000 0.000 63.000 88.700 ;
        RECT  0.600 0.600 1.480 91.220 ;
        RECT  0.600 90.750 64.400 91.220 ;
        LAYER TOP_M ;
        RECT  0.600 247.690 64.400 248.850 ;
        RECT  0.600 247.690 23.010 249.400 ;
        RECT  26.470 247.690 27.110 249.400 ;
        RECT  30.330 247.690 64.400 249.400 ;
        RECT  2.000 0.000 63.000 91.190 ;
        RECT  0.600 0.600 64.400 91.190 ;
    END
END pc3t01d

MACRO pc3t01
    CLASS PAD ;
    FOREIGN pc3t01 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 65.000 BY 250.000 ;
    SYMMETRY X Y R90 ;
    SITE IOSite_c ;
    PIN PAD
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 55.440  LAYER TOP_M  ;
        ANTENNAPARTIALMETALSIDEAREA 287.938  LAYER M3  ;
        ANTENNAPARTIALMETALSIDEAREA 480.740  LAYER M2  ;
        ANTENNADIFFAREA 2657.280  LAYER TOP_M  ;
        ANTENNADIFFAREA 2657.280  LAYER M3  ;
        ANTENNADIFFAREA 1209.600  LAYER M2  ;
        ANTENNAPARTIALCUTAREA 632.318  LAYER TOP_V  ;
        ANTENNAPARTIALCUTAREA 349.898  LAYER V3  ;
        ANTENNAPARTIALCUTAREA 255.798  LAYER V2  ;
        PORT
        LAYER M3 ;
        RECT  23.740 249.580 25.740 250.000 ;
        LAYER M2 ;
        RECT  2.000 61.000 63.000 90.230 ;
        RECT  23.740 246.275 25.740 250.000 ;
        END
    END PAD
    PIN OEN
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 81.726  LAYER M2  ;
        ANTENNAPARTIALMETALSIDEAREA 67.374  LAYER M1  ;
        ANTENNAPARTIALMETALSIDEAREA 41.679  LAYER M3  ;
        ANTENNADIFFAREA 0.250  LAYER M3  ;
        ANTENNAPARTIALCUTAREA 0.135  LAYER V3  ;
        ANTENNAPARTIALCUTAREA 0.203  LAYER V2  ;
        ANTENNAGATEAREA 8.100  LAYER M2  ;
        ANTENNAGATEAREA 9.900  LAYER M3  ;
        PORT
        LAYER M3 ;
        RECT  28.870 249.580 29.600 250.000 ;
        LAYER M2 ;
        RECT  28.870 249.580 29.600 250.000 ;
        END
    END OEN
    PIN I
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 80.804  LAYER M2  ;
        ANTENNAPARTIALMETALSIDEAREA 67.374  LAYER M1  ;
        ANTENNAPARTIALMETALSIDEAREA 41.096  LAYER M3  ;
        ANTENNADIFFAREA 0.250  LAYER M3  ;
        ANTENNAPARTIALCUTAREA 0.135  LAYER V3  ;
        ANTENNAPARTIALCUTAREA 0.203  LAYER V2  ;
        ANTENNAGATEAREA 8.100  LAYER M2  ;
        ANTENNAGATEAREA 9.900  LAYER M3  ;
        PORT
        LAYER M3 ;
        RECT  27.840 249.580 28.570 250.000 ;
        LAYER M2 ;
        RECT  27.840 249.580 28.570 250.000 ;
        END
    END I
    PIN VDDO
        DIRECTION INOUT ;
        USE power ;
        PORT
        LAYER M3 ;
        RECT  64.200 192.330 65.000 200.640 ;
        RECT  0.000 201.660 65.000 221.520 ;
        RECT  0.000 222.720 65.000 246.820 ;
        RECT  0.000 192.330 0.800 200.640 ;
        LAYER M2 ;
        RECT  0.000 186.470 65.000 195.650 ;
        LAYER TOP_M ;
        RECT  0.000 195.170 65.000 200.640 ;
        RECT  0.000 201.660 65.000 221.520 ;
        RECT  0.000 222.720 65.000 246.820 ;
        END
    END VDDO
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        PORT
        LAYER M3 ;
        RECT  64.200 163.510 65.000 190.890 ;
        RECT  0.000 163.510 0.800 190.890 ;
        LAYER M2 ;
        RECT  0.000 172.080 65.000 183.060 ;
        LAYER TOP_M ;
        RECT  0.000 163.500 65.000 194.560 ;
        END
    END VDD
    PIN VSSO
        DIRECTION INOUT ;
        USE ground ;
        PORT
        LAYER M3 ;
        RECT  0.000 92.060 65.000 123.250 ;
        RECT  64.200 149.940 65.000 162.610 ;
        RECT  0.000 149.940 0.800 162.610 ;
        LAYER M2 ;
        RECT  0.000 147.040 65.000 154.520 ;
        LAYER TOP_M ;
        RECT  0.000 92.060 65.000 123.250 ;
        RECT  0.000 155.410 65.000 162.610 ;
        END
    END VSSO
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        PORT
        LAYER M3 ;
        RECT  64.200 130.690 65.000 148.880 ;
        RECT  0.000 130.690 0.800 148.880 ;
        LAYER M2 ;
        RECT  0.000 136.310 65.000 146.340 ;
        LAYER TOP_M ;
        RECT  0.000 123.850 65.000 154.560 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  2.000 0.000 63.000 250.000 ;
        RECT  0.000 88.990 65.000 130.360 ;
        RECT  0.000 136.510 65.000 157.550 ;
        RECT  0.315 158.150 64.700 158.460 ;
        RECT  0.300 158.930 64.700 159.230 ;
        RECT  0.300 159.530 64.700 159.830 ;
        RECT  0.300 160.130 64.700 160.430 ;
        RECT  0.300 160.730 64.700 161.030 ;
        RECT  0.300 161.330 64.700 161.630 ;
        RECT  0.300 161.910 64.700 162.190 ;
        RECT  0.300 162.490 64.700 162.770 ;
        RECT  0.300 163.070 64.700 163.350 ;
        RECT  0.300 163.650 64.700 163.950 ;
        RECT  0.300 164.250 64.700 164.550 ;
        RECT  0.300 164.850 64.700 165.150 ;
        RECT  0.300 165.450 64.700 165.750 ;
        RECT  0.300 166.050 64.700 166.350 ;
        RECT  0.300 166.650 64.700 166.960 ;
        RECT  0.300 167.260 64.700 167.560 ;
        RECT  0.300 167.860 64.700 168.160 ;
        RECT  0.000 169.150 65.000 197.240 ;
        RECT  0.600 0.600 64.400 250.000 ;
        RECT  0.000 198.470 65.000 250.000 ;
        LAYER M2 ;
        RECT  63.180 196.430 63.670 249.400 ;
        RECT  0.600 196.440 64.400 245.485 ;
        RECT  26.530 196.440 64.400 248.790 ;
        RECT  0.600 196.440 22.950 249.400 ;
        RECT  26.530 196.440 27.050 249.400 ;
        RECT  30.390 196.440 64.400 249.400 ;
        RECT  0.600 183.850 64.400 185.680 ;
        RECT  46.230 183.850 51.730 185.870 ;
        RECT  19.790 155.160 20.140 171.290 ;
        RECT  20.440 155.140 20.760 171.290 ;
        RECT  53.655 155.035 53.935 171.290 ;
        RECT  56.365 155.280 56.645 171.290 ;
        RECT  57.120 155.300 57.400 171.290 ;
        RECT  57.835 155.130 58.115 171.290 ;
        RECT  0.600 155.310 64.400 171.290 ;
        RECT  53.895 155.310 55.870 171.370 ;
        RECT  3.210 155.310 3.490 171.380 ;
        RECT  34.655 155.310 38.715 171.480 ;
        RECT  39.605 155.310 42.020 171.480 ;
        RECT  2.000 0.000 63.000 60.210 ;
        RECT  0.600 0.600 64.400 60.210 ;
        RECT  0.600 0.600 1.210 135.520 ;
        RECT  0.600 91.020 64.400 135.520 ;
        RECT  4.080 91.020 60.940 135.690 ;
        RECT  62.580 91.020 62.995 135.710 ;
        LAYER M3 ;
        RECT  0.600 247.660 23.220 248.740 ;
        RECT  0.600 247.660 22.900 249.400 ;
        RECT  26.260 247.660 64.400 248.740 ;
        RECT  26.580 247.660 27.000 249.400 ;
        RECT  30.440 247.660 64.400 249.400 ;
        RECT  0.600 124.090 64.400 129.850 ;
        RECT  3.990 123.970 60.900 135.790 ;
        RECT  1.640 124.090 63.600 135.790 ;
        RECT  1.810 124.090 2.830 154.520 ;
        RECT  5.155 123.970 60.900 171.560 ;
        RECT  1.640 155.040 63.600 171.560 ;
        RECT  1.640 183.580 63.600 185.950 ;
        RECT  5.490 124.090 63.600 200.820 ;
        RECT  1.640 196.170 63.600 200.820 ;
        RECT  0.600 0.600 64.400 60.480 ;
        RECT  2.000 0.000 63.000 88.700 ;
        RECT  0.600 0.600 1.480 91.220 ;
        RECT  0.600 90.750 64.400 91.220 ;
        LAYER TOP_M ;
        RECT  0.600 247.690 64.400 248.850 ;
        RECT  0.600 247.690 23.010 249.400 ;
        RECT  26.470 247.690 27.110 249.400 ;
        RECT  30.330 247.690 64.400 249.400 ;
        RECT  2.000 0.000 63.000 91.190 ;
        RECT  0.600 0.600 64.400 91.190 ;
    END
END pc3t01

MACRO pc3o05
    CLASS PAD ;
    FOREIGN pc3o05 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 65.000 BY 250.000 ;
    SYMMETRY X Y R90 ;
    SITE IOSite_c ;
    PIN PAD
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 55.440  LAYER TOP_M  ;
        ANTENNAPARTIALMETALSIDEAREA 287.938  LAYER M3  ;
        ANTENNAPARTIALMETALSIDEAREA 480.740  LAYER M2  ;
        ANTENNADIFFAREA 2657.280  LAYER TOP_M  ;
        ANTENNADIFFAREA 2657.280  LAYER M3  ;
        ANTENNADIFFAREA 1209.600  LAYER M2  ;
        ANTENNAPARTIALCUTAREA 632.318  LAYER TOP_V  ;
        ANTENNAPARTIALCUTAREA 349.898  LAYER V3  ;
        ANTENNAPARTIALCUTAREA 255.798  LAYER V2  ;
        PORT
        LAYER M3 ;
        RECT  26.310 249.580 28.310 250.000 ;
        LAYER M2 ;
        RECT  2.000 61.000 63.000 90.230 ;
        RECT  26.310 246.275 28.310 250.000 ;
        END
    END PAD
    PIN I
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 67.374  LAYER M1  ;
        ANTENNAPARTIALMETALSIDEAREA 81.652  LAYER M2  ;
        ANTENNAPARTIALMETALSIDEAREA 41.425  LAYER M3  ;
        ANTENNADIFFAREA 0.250  LAYER M3  ;
        ANTENNAPARTIALCUTAREA 0.338  LAYER V2  ;
        ANTENNAPARTIALCUTAREA 0.135  LAYER V3  ;
        ANTENNAGATEAREA 18.900  LAYER M2  ;
        ANTENNAGATEAREA 20.700  LAYER M3  ;
        PORT
        LAYER M3 ;
        RECT  30.310 249.580 31.040 250.000 ;
        LAYER M2 ;
        RECT  30.310 249.580 31.040 250.000 ;
        END
    END I
    PIN VDDO
        DIRECTION INOUT ;
        USE power ;
        PORT
        LAYER M3 ;
        RECT  64.200 192.330 65.000 200.640 ;
        RECT  0.000 201.660 65.000 221.520 ;
        RECT  0.000 222.720 65.000 246.820 ;
        RECT  0.000 192.330 0.800 200.640 ;
        LAYER M2 ;
        RECT  0.000 186.470 65.000 195.650 ;
        LAYER TOP_M ;
        RECT  0.000 195.170 65.000 200.640 ;
        RECT  0.000 201.660 65.000 221.520 ;
        RECT  0.000 222.720 65.000 246.820 ;
        END
    END VDDO
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        PORT
        LAYER M3 ;
        RECT  64.200 163.510 65.000 190.890 ;
        RECT  0.000 163.510 0.800 190.890 ;
        LAYER M2 ;
        RECT  0.000 172.080 65.000 183.060 ;
        LAYER TOP_M ;
        RECT  0.000 163.500 65.000 194.560 ;
        END
    END VDD
    PIN VSSO
        DIRECTION INOUT ;
        USE ground ;
        PORT
        LAYER M3 ;
        RECT  0.000 92.060 65.000 123.250 ;
        RECT  64.200 149.940 65.000 162.610 ;
        RECT  0.000 149.940 0.800 162.610 ;
        LAYER M2 ;
        RECT  0.000 147.040 65.000 154.520 ;
        LAYER TOP_M ;
        RECT  0.000 92.060 65.000 123.250 ;
        RECT  0.000 155.410 65.000 162.610 ;
        END
    END VSSO
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        PORT
        LAYER M3 ;
        RECT  64.200 130.690 65.000 148.880 ;
        RECT  0.000 130.690 0.800 148.880 ;
        LAYER M2 ;
        RECT  0.000 136.310 65.000 146.340 ;
        LAYER TOP_M ;
        RECT  0.000 123.850 65.000 154.560 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  2.000 0.000 63.000 250.000 ;
        RECT  0.000 88.990 65.000 130.360 ;
        RECT  0.000 136.510 65.000 157.550 ;
        RECT  0.300 158.930 64.700 159.230 ;
        RECT  0.300 159.530 64.700 159.830 ;
        RECT  0.300 160.130 64.700 160.430 ;
        RECT  0.300 160.730 64.700 161.030 ;
        RECT  0.300 161.330 64.700 161.630 ;
        RECT  0.300 161.910 64.700 162.190 ;
        RECT  0.300 162.490 64.700 162.770 ;
        RECT  0.300 163.070 64.700 163.350 ;
        RECT  0.300 163.650 64.700 163.950 ;
        RECT  0.300 164.250 64.700 164.550 ;
        RECT  0.300 164.850 64.700 165.150 ;
        RECT  0.300 165.450 64.700 165.750 ;
        RECT  0.300 166.050 64.700 166.350 ;
        RECT  0.300 166.650 64.700 166.960 ;
        RECT  0.300 167.260 64.700 167.560 ;
        RECT  0.300 167.860 64.700 168.160 ;
        RECT  0.000 169.150 65.000 197.240 ;
        RECT  0.600 0.600 64.400 250.000 ;
        RECT  0.000 198.470 65.000 250.000 ;
        LAYER M2 ;
        RECT  2.800 196.110 3.220 249.400 ;
        RECT  63.180 196.430 63.670 249.400 ;
        RECT  0.600 196.440 64.400 245.485 ;
        RECT  29.100 196.440 64.400 248.790 ;
        RECT  0.600 196.440 25.520 249.400 ;
        RECT  29.100 196.440 29.520 249.400 ;
        RECT  31.830 196.440 64.400 249.400 ;
        RECT  55.890 183.790 56.190 185.680 ;
        RECT  58.060 183.750 58.350 185.680 ;
        RECT  0.600 183.850 64.400 185.680 ;
        RECT  46.070 183.850 51.600 185.820 ;
        RECT  8.170 155.125 8.490 171.290 ;
        RECT  43.245 155.035 43.525 171.290 ;
        RECT  45.955 155.280 46.235 171.370 ;
        RECT  47.425 155.130 47.705 171.370 ;
        RECT  58.295 155.175 58.605 171.290 ;
        RECT  60.755 155.175 61.065 171.290 ;
        RECT  63.290 155.270 63.600 171.290 ;
        RECT  0.600 155.310 64.400 171.290 ;
        RECT  43.485 155.310 56.355 171.370 ;
        RECT  29.195 155.310 31.610 171.480 ;
        RECT  2.000 0.000 63.000 60.210 ;
        RECT  0.600 0.600 64.400 60.210 ;
        RECT  0.600 0.600 1.210 135.520 ;
        RECT  0.600 91.020 64.400 135.520 ;
        RECT  4.080 91.020 60.940 135.690 ;
        LAYER M3 ;
        RECT  0.600 247.660 25.790 248.740 ;
        RECT  0.600 247.660 25.470 249.400 ;
        RECT  28.830 247.660 64.400 248.740 ;
        RECT  29.150 247.660 29.470 249.400 ;
        RECT  31.880 247.660 64.400 249.400 ;
        RECT  4.040 123.850 60.900 200.820 ;
        RECT  0.600 124.090 64.400 129.850 ;
        RECT  1.640 124.090 63.600 135.790 ;
        RECT  1.810 124.090 2.830 154.520 ;
        RECT  1.640 155.040 63.600 171.560 ;
        RECT  1.640 183.580 63.600 185.950 ;
        RECT  2.800 155.040 63.600 200.820 ;
        RECT  3.340 124.090 63.600 200.820 ;
        RECT  1.640 196.170 63.600 200.820 ;
        RECT  0.600 0.600 64.400 60.480 ;
        RECT  2.000 0.000 63.000 88.700 ;
        RECT  0.600 0.600 1.480 91.220 ;
        RECT  0.600 90.750 64.400 91.220 ;
        LAYER TOP_M ;
        RECT  0.600 247.690 64.400 248.850 ;
        RECT  0.600 247.690 25.580 249.400 ;
        RECT  29.040 247.690 29.580 249.400 ;
        RECT  31.770 247.690 64.400 249.400 ;
        RECT  2.000 0.000 63.000 91.190 ;
        RECT  0.600 0.600 64.400 91.190 ;
    END
END pc3o05

MACRO pc3o04
    CLASS PAD ;
    FOREIGN pc3o04 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 65.000 BY 250.000 ;
    SYMMETRY X Y R90 ;
    SITE IOSite_c ;
    PIN PAD
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 55.440  LAYER TOP_M  ;
        ANTENNAPARTIALMETALSIDEAREA 287.938  LAYER M3  ;
        ANTENNAPARTIALMETALSIDEAREA 480.740  LAYER M2  ;
        ANTENNADIFFAREA 2657.280  LAYER TOP_M  ;
        ANTENNADIFFAREA 2657.280  LAYER M3  ;
        ANTENNADIFFAREA 1209.600  LAYER M2  ;
        ANTENNAPARTIALCUTAREA 632.318  LAYER TOP_V  ;
        ANTENNAPARTIALCUTAREA 349.898  LAYER V3  ;
        ANTENNAPARTIALCUTAREA 255.798  LAYER V2  ;
        PORT
        LAYER M3 ;
        RECT  26.310 249.580 28.310 250.000 ;
        LAYER M2 ;
        RECT  2.000 61.000 63.000 90.230 ;
        RECT  26.310 246.275 28.310 250.000 ;
        END
    END PAD
    PIN I
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 67.374  LAYER M1  ;
        ANTENNAPARTIALMETALSIDEAREA 81.652  LAYER M2  ;
        ANTENNAPARTIALMETALSIDEAREA 41.425  LAYER M3  ;
        ANTENNADIFFAREA 0.250  LAYER M3  ;
        ANTENNAPARTIALCUTAREA 0.338  LAYER V2  ;
        ANTENNAPARTIALCUTAREA 0.135  LAYER V3  ;
        ANTENNAGATEAREA 18.900  LAYER M2  ;
        ANTENNAGATEAREA 20.700  LAYER M3  ;
        PORT
        LAYER M3 ;
        RECT  30.310 249.580 31.040 250.000 ;
        LAYER M2 ;
        RECT  30.310 249.580 31.040 250.000 ;
        END
    END I
    PIN VDDO
        DIRECTION INOUT ;
        USE power ;
        PORT
        LAYER M3 ;
        RECT  64.200 192.330 65.000 200.640 ;
        RECT  0.000 201.660 65.000 221.520 ;
        RECT  0.000 222.720 65.000 246.820 ;
        RECT  0.000 192.330 0.800 200.640 ;
        LAYER M2 ;
        RECT  0.000 186.470 65.000 195.650 ;
        LAYER TOP_M ;
        RECT  0.000 195.170 65.000 200.640 ;
        RECT  0.000 201.660 65.000 221.520 ;
        RECT  0.000 222.720 65.000 246.820 ;
        END
    END VDDO
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        PORT
        LAYER M3 ;
        RECT  64.200 163.510 65.000 190.890 ;
        RECT  0.000 163.510 0.800 190.890 ;
        LAYER M2 ;
        RECT  0.000 172.080 65.000 183.060 ;
        LAYER TOP_M ;
        RECT  0.000 163.500 65.000 194.560 ;
        END
    END VDD
    PIN VSSO
        DIRECTION INOUT ;
        USE ground ;
        PORT
        LAYER M3 ;
        RECT  0.000 92.060 65.000 123.250 ;
        RECT  64.200 149.940 65.000 162.610 ;
        RECT  0.000 149.940 0.800 162.610 ;
        LAYER M2 ;
        RECT  0.000 147.040 65.000 154.520 ;
        LAYER TOP_M ;
        RECT  0.000 92.060 65.000 123.250 ;
        RECT  0.000 155.410 65.000 162.610 ;
        END
    END VSSO
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        PORT
        LAYER M3 ;
        RECT  64.200 130.690 65.000 148.880 ;
        RECT  0.000 130.690 0.800 148.880 ;
        LAYER M2 ;
        RECT  0.000 136.310 65.000 146.340 ;
        LAYER TOP_M ;
        RECT  0.000 123.850 65.000 154.560 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  2.000 0.000 63.000 250.000 ;
        RECT  0.000 88.990 65.000 130.360 ;
        RECT  0.000 136.510 65.000 157.550 ;
        RECT  0.300 158.930 64.700 159.230 ;
        RECT  0.300 159.530 64.700 159.830 ;
        RECT  0.300 160.130 64.700 160.430 ;
        RECT  0.300 160.730 64.700 161.030 ;
        RECT  0.300 161.330 64.700 161.630 ;
        RECT  0.300 161.910 64.700 162.190 ;
        RECT  0.300 162.490 64.700 162.770 ;
        RECT  0.300 163.070 64.700 163.350 ;
        RECT  0.300 163.650 64.700 163.950 ;
        RECT  0.300 164.250 64.700 164.550 ;
        RECT  0.300 164.850 64.700 165.150 ;
        RECT  0.300 165.450 64.700 165.750 ;
        RECT  0.300 166.050 64.700 166.350 ;
        RECT  0.300 166.650 64.700 166.960 ;
        RECT  0.300 167.260 64.700 167.560 ;
        RECT  0.300 167.860 64.700 168.160 ;
        RECT  0.000 169.150 65.000 197.240 ;
        RECT  0.600 0.600 64.400 250.000 ;
        RECT  0.000 198.470 65.000 250.000 ;
        LAYER M2 ;
        RECT  63.180 196.430 63.670 249.400 ;
        RECT  0.600 196.440 64.400 245.485 ;
        RECT  29.100 196.440 64.400 248.790 ;
        RECT  0.600 196.440 25.520 249.400 ;
        RECT  29.100 196.440 29.520 249.400 ;
        RECT  31.830 196.440 64.400 249.400 ;
        RECT  55.890 183.790 56.190 185.680 ;
        RECT  58.060 183.750 58.350 185.680 ;
        RECT  0.600 183.850 64.400 185.680 ;
        RECT  46.070 183.850 51.600 185.820 ;
        RECT  8.170 155.125 8.490 171.290 ;
        RECT  43.245 155.035 43.525 171.290 ;
        RECT  45.955 155.280 46.235 171.370 ;
        RECT  47.425 155.130 47.705 171.370 ;
        RECT  58.165 155.175 58.475 171.290 ;
        RECT  60.625 155.175 60.935 171.290 ;
        RECT  63.160 155.270 63.470 171.290 ;
        RECT  0.600 155.310 64.400 171.290 ;
        RECT  43.485 155.310 56.355 171.370 ;
        RECT  29.195 155.310 31.610 171.480 ;
        RECT  2.000 0.000 63.000 60.210 ;
        RECT  0.600 0.600 64.400 60.210 ;
        RECT  0.600 0.600 1.210 135.520 ;
        RECT  0.600 91.020 64.400 135.520 ;
        RECT  4.080 91.020 60.940 135.690 ;
        LAYER M3 ;
        RECT  0.600 247.660 25.790 248.740 ;
        RECT  0.600 247.660 25.470 249.400 ;
        RECT  28.830 247.660 64.400 248.740 ;
        RECT  29.150 247.660 29.470 249.400 ;
        RECT  31.880 247.660 64.400 249.400 ;
        RECT  0.600 124.090 64.400 129.850 ;
        RECT  1.640 124.090 63.600 135.790 ;
        RECT  1.810 124.090 2.830 154.520 ;
        RECT  1.640 155.040 63.600 171.560 ;
        RECT  1.640 183.580 63.600 185.950 ;
        RECT  2.800 155.040 63.600 200.820 ;
        RECT  3.215 124.090 63.600 200.820 ;
        RECT  1.640 196.170 63.600 200.820 ;
        RECT  0.600 0.600 64.400 60.480 ;
        RECT  2.000 0.000 63.000 88.700 ;
        RECT  0.600 0.600 1.480 91.220 ;
        RECT  0.600 90.750 64.400 91.220 ;
        LAYER TOP_M ;
        RECT  0.600 247.690 64.400 248.850 ;
        RECT  0.600 247.690 25.580 249.400 ;
        RECT  29.040 247.690 29.580 249.400 ;
        RECT  31.770 247.690 64.400 249.400 ;
        RECT  2.000 0.000 63.000 91.190 ;
        RECT  0.600 0.600 64.400 91.190 ;
    END
END pc3o04

MACRO pc3o03
    CLASS PAD ;
    FOREIGN pc3o03 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 65.000 BY 250.000 ;
    SYMMETRY X Y R90 ;
    SITE IOSite_c ;
    PIN PAD
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 55.440  LAYER TOP_M  ;
        ANTENNAPARTIALMETALSIDEAREA 287.938  LAYER M3  ;
        ANTENNAPARTIALMETALSIDEAREA 480.740  LAYER M2  ;
        ANTENNADIFFAREA 2657.280  LAYER TOP_M  ;
        ANTENNADIFFAREA 2657.280  LAYER M3  ;
        ANTENNADIFFAREA 1209.600  LAYER M2  ;
        ANTENNAPARTIALCUTAREA 632.318  LAYER TOP_V  ;
        ANTENNAPARTIALCUTAREA 349.898  LAYER V3  ;
        ANTENNAPARTIALCUTAREA 255.798  LAYER V2  ;
        PORT
        LAYER M3 ;
        RECT  26.310 249.580 28.310 250.000 ;
        LAYER M2 ;
        RECT  2.000 61.000 63.000 90.230 ;
        RECT  26.310 246.275 28.310 250.000 ;
        END
    END PAD
    PIN I
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 67.374  LAYER M1  ;
        ANTENNAPARTIALMETALSIDEAREA 81.652  LAYER M2  ;
        ANTENNAPARTIALMETALSIDEAREA 41.425  LAYER M3  ;
        ANTENNADIFFAREA 0.250  LAYER M3  ;
        ANTENNAPARTIALCUTAREA 0.338  LAYER V2  ;
        ANTENNAPARTIALCUTAREA 0.135  LAYER V3  ;
        ANTENNAGATEAREA 18.900  LAYER M2  ;
        ANTENNAGATEAREA 20.700  LAYER M3  ;
        PORT
        LAYER M3 ;
        RECT  30.310 249.580 31.040 250.000 ;
        LAYER M2 ;
        RECT  30.310 249.580 31.040 250.000 ;
        END
    END I
    PIN VDDO
        DIRECTION INOUT ;
        USE power ;
        PORT
        LAYER M3 ;
        RECT  64.200 192.330 65.000 200.640 ;
        RECT  0.000 201.660 65.000 221.520 ;
        RECT  0.000 222.720 65.000 246.820 ;
        RECT  0.000 192.330 0.800 200.640 ;
        LAYER M2 ;
        RECT  0.000 186.470 65.000 195.650 ;
        LAYER TOP_M ;
        RECT  0.000 195.170 65.000 200.640 ;
        RECT  0.000 201.660 65.000 221.520 ;
        RECT  0.000 222.720 65.000 246.820 ;
        END
    END VDDO
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        PORT
        LAYER M3 ;
        RECT  64.200 163.510 65.000 190.890 ;
        RECT  0.000 163.510 0.800 190.890 ;
        LAYER M2 ;
        RECT  0.000 172.080 65.000 183.060 ;
        LAYER TOP_M ;
        RECT  0.000 163.500 65.000 194.560 ;
        END
    END VDD
    PIN VSSO
        DIRECTION INOUT ;
        USE ground ;
        PORT
        LAYER M3 ;
        RECT  0.000 92.060 65.000 123.250 ;
        RECT  64.200 149.940 65.000 162.610 ;
        RECT  0.000 149.940 0.800 162.610 ;
        LAYER M2 ;
        RECT  0.000 147.040 65.000 154.520 ;
        LAYER TOP_M ;
        RECT  0.000 92.060 65.000 123.250 ;
        RECT  0.000 155.410 65.000 162.610 ;
        END
    END VSSO
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        PORT
        LAYER M3 ;
        RECT  64.200 130.690 65.000 148.880 ;
        RECT  0.000 130.690 0.800 148.880 ;
        LAYER M2 ;
        RECT  0.000 136.310 65.000 146.340 ;
        LAYER TOP_M ;
        RECT  0.000 123.850 65.000 154.560 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  2.000 0.000 63.000 250.000 ;
        RECT  0.000 88.990 65.000 130.360 ;
        RECT  0.000 136.510 65.000 157.550 ;
        RECT  0.300 158.930 64.700 159.230 ;
        RECT  0.300 159.530 64.700 159.830 ;
        RECT  0.300 160.130 64.700 160.430 ;
        RECT  0.300 160.730 64.700 161.030 ;
        RECT  0.300 161.330 64.700 161.630 ;
        RECT  0.300 161.910 64.700 162.190 ;
        RECT  0.300 162.490 64.700 162.770 ;
        RECT  0.300 163.070 64.700 163.350 ;
        RECT  0.300 163.650 64.700 163.950 ;
        RECT  0.300 164.250 64.700 164.550 ;
        RECT  0.300 164.850 64.700 165.150 ;
        RECT  0.300 165.450 64.700 165.750 ;
        RECT  0.300 166.050 64.700 166.350 ;
        RECT  0.300 166.650 64.700 166.960 ;
        RECT  0.300 167.260 64.700 167.560 ;
        RECT  0.300 167.860 64.700 168.160 ;
        RECT  0.000 169.150 65.000 197.240 ;
        RECT  0.600 0.600 64.400 250.000 ;
        RECT  0.000 198.470 65.000 250.000 ;
        LAYER M2 ;
        RECT  2.800 196.110 3.220 249.400 ;
        RECT  63.180 196.430 63.670 249.400 ;
        RECT  0.600 196.440 64.400 245.485 ;
        RECT  29.100 196.440 64.400 248.790 ;
        RECT  0.600 196.440 25.520 249.400 ;
        RECT  29.100 196.440 29.520 249.400 ;
        RECT  31.830 196.440 64.400 249.400 ;
        RECT  55.890 183.790 56.190 185.680 ;
        RECT  58.060 183.750 58.350 185.680 ;
        RECT  0.600 183.850 64.400 185.680 ;
        RECT  46.070 183.850 51.600 185.820 ;
        RECT  8.170 155.125 8.490 171.290 ;
        RECT  43.245 155.035 43.525 171.290 ;
        RECT  45.955 155.280 46.235 171.370 ;
        RECT  47.425 155.130 47.705 171.370 ;
        RECT  58.045 155.175 58.355 171.290 ;
        RECT  60.505 155.175 60.815 171.290 ;
        RECT  63.040 155.270 63.350 171.290 ;
        RECT  0.600 155.310 64.400 171.290 ;
        RECT  43.485 155.310 56.355 171.370 ;
        RECT  29.195 155.310 31.610 171.480 ;
        RECT  2.000 0.000 63.000 60.210 ;
        RECT  0.600 0.600 64.400 60.210 ;
        RECT  0.600 0.600 1.210 135.520 ;
        RECT  0.600 91.020 64.400 135.520 ;
        RECT  4.080 91.020 60.940 135.690 ;
        LAYER M3 ;
        RECT  0.600 247.660 25.790 248.740 ;
        RECT  0.600 247.660 25.470 249.400 ;
        RECT  28.830 247.660 64.400 248.740 ;
        RECT  29.150 247.660 29.470 249.400 ;
        RECT  31.880 247.660 64.400 249.400 ;
        RECT  4.040 123.970 60.900 200.820 ;
        RECT  0.600 124.090 64.400 129.850 ;
        RECT  1.640 124.090 63.600 135.790 ;
        RECT  1.810 124.090 2.830 154.520 ;
        RECT  1.640 155.040 63.600 171.560 ;
        RECT  1.640 183.580 63.600 185.950 ;
        RECT  2.800 155.040 63.600 200.820 ;
        RECT  3.230 124.090 63.600 200.820 ;
        RECT  1.640 196.170 63.600 200.820 ;
        RECT  0.600 0.600 64.400 60.480 ;
        RECT  2.000 0.000 63.000 88.700 ;
        RECT  0.600 0.600 1.480 91.220 ;
        RECT  0.600 90.750 64.400 91.220 ;
        LAYER TOP_M ;
        RECT  0.600 247.690 64.400 248.850 ;
        RECT  0.600 247.690 25.580 249.400 ;
        RECT  29.040 247.690 29.580 249.400 ;
        RECT  31.770 247.690 64.400 249.400 ;
        RECT  2.000 0.000 63.000 91.190 ;
        RECT  0.600 0.600 64.400 91.190 ;
    END
END pc3o03

MACRO pc3o02
    CLASS PAD ;
    FOREIGN pc3o02 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 65.000 BY 250.000 ;
    SYMMETRY X Y R90 ;
    SITE IOSite_c ;
    PIN PAD
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 55.440  LAYER TOP_M  ;
        ANTENNAPARTIALMETALSIDEAREA 287.938  LAYER M3  ;
        ANTENNAPARTIALMETALSIDEAREA 480.740  LAYER M2  ;
        ANTENNADIFFAREA 2657.280  LAYER TOP_M  ;
        ANTENNADIFFAREA 2657.280  LAYER M3  ;
        ANTENNADIFFAREA 1209.600  LAYER M2  ;
        ANTENNAPARTIALCUTAREA 632.318  LAYER TOP_V  ;
        ANTENNAPARTIALCUTAREA 349.898  LAYER V3  ;
        ANTENNAPARTIALCUTAREA 255.798  LAYER V2  ;
        PORT
        LAYER M3 ;
        RECT  26.310 249.580 28.310 250.000 ;
        LAYER M2 ;
        RECT  2.000 61.000 63.000 90.230 ;
        RECT  26.310 246.275 28.310 250.000 ;
        END
    END PAD
    PIN I
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 67.374  LAYER M1  ;
        ANTENNAPARTIALMETALSIDEAREA 81.652  LAYER M2  ;
        ANTENNAPARTIALMETALSIDEAREA 41.425  LAYER M3  ;
        ANTENNADIFFAREA 0.250  LAYER M3  ;
        ANTENNAPARTIALCUTAREA 0.135  LAYER V3  ;
        ANTENNAPARTIALCUTAREA 0.338  LAYER V2  ;
        ANTENNAGATEAREA 18.900  LAYER M2  ;
        ANTENNAGATEAREA 20.700  LAYER M3  ;
        PORT
        LAYER M3 ;
        RECT  30.310 249.580 31.040 250.000 ;
        LAYER M2 ;
        RECT  30.310 249.580 31.040 250.000 ;
        END
    END I
    PIN VDDO
        DIRECTION INOUT ;
        USE power ;
        PORT
        LAYER M3 ;
        RECT  64.200 192.330 65.000 200.640 ;
        RECT  0.000 201.660 65.000 221.520 ;
        RECT  0.000 222.720 65.000 246.820 ;
        RECT  0.000 192.330 0.800 200.640 ;
        LAYER M2 ;
        RECT  0.000 186.470 65.000 195.650 ;
        LAYER TOP_M ;
        RECT  0.000 195.170 65.000 200.640 ;
        RECT  0.000 201.660 65.000 221.520 ;
        RECT  0.000 222.720 65.000 246.820 ;
        END
    END VDDO
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        PORT
        LAYER M3 ;
        RECT  64.200 163.510 65.000 190.890 ;
        RECT  0.000 163.510 0.800 190.890 ;
        LAYER M2 ;
        RECT  0.000 172.080 65.000 183.060 ;
        LAYER TOP_M ;
        RECT  0.000 163.500 65.000 194.560 ;
        END
    END VDD
    PIN VSSO
        DIRECTION INOUT ;
        USE ground ;
        PORT
        LAYER M3 ;
        RECT  0.000 92.060 65.000 123.250 ;
        RECT  64.200 149.940 65.000 162.610 ;
        RECT  0.000 149.940 0.800 162.610 ;
        LAYER M2 ;
        RECT  0.000 147.040 65.000 154.520 ;
        LAYER TOP_M ;
        RECT  0.000 92.060 65.000 123.250 ;
        RECT  0.000 155.410 65.000 162.610 ;
        END
    END VSSO
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        PORT
        LAYER M3 ;
        RECT  64.200 130.690 65.000 148.880 ;
        RECT  0.000 130.690 0.800 148.880 ;
        LAYER M2 ;
        RECT  0.000 136.310 65.000 146.340 ;
        LAYER TOP_M ;
        RECT  0.000 123.850 65.000 154.560 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  2.000 0.000 63.000 250.000 ;
        RECT  0.000 88.990 65.000 130.360 ;
        RECT  0.000 136.510 65.000 157.550 ;
        RECT  0.300 158.930 64.700 159.230 ;
        RECT  0.300 159.530 64.700 159.830 ;
        RECT  0.300 160.130 64.700 160.430 ;
        RECT  0.300 160.730 64.700 161.030 ;
        RECT  0.300 161.330 64.700 161.630 ;
        RECT  0.300 161.910 64.700 162.190 ;
        RECT  0.300 162.490 64.700 162.770 ;
        RECT  0.300 163.070 64.700 163.350 ;
        RECT  0.300 163.650 64.700 163.950 ;
        RECT  0.300 164.250 64.700 164.550 ;
        RECT  0.300 164.850 64.700 165.150 ;
        RECT  0.300 165.450 64.700 165.750 ;
        RECT  0.300 166.050 64.700 166.350 ;
        RECT  0.300 166.650 64.700 166.960 ;
        RECT  0.300 167.260 64.700 167.560 ;
        RECT  0.300 167.860 64.700 168.160 ;
        RECT  0.000 169.150 65.000 197.240 ;
        RECT  0.600 0.600 64.400 250.000 ;
        RECT  0.000 198.470 65.000 250.000 ;
        LAYER M2 ;
        RECT  2.790 196.270 3.210 249.400 ;
        RECT  63.180 196.430 63.670 249.400 ;
        RECT  0.600 196.440 64.400 245.485 ;
        RECT  29.100 196.440 64.400 248.790 ;
        RECT  0.600 196.440 25.520 249.400 ;
        RECT  29.100 196.440 29.520 249.400 ;
        RECT  31.830 196.440 64.400 249.400 ;
        RECT  55.890 183.790 56.190 185.680 ;
        RECT  58.060 183.750 58.350 185.680 ;
        RECT  0.600 183.850 64.400 185.680 ;
        RECT  46.070 183.850 51.600 185.820 ;
        RECT  7.575 155.125 7.895 171.290 ;
        RECT  43.245 155.035 43.525 171.290 ;
        RECT  45.955 155.280 46.235 171.370 ;
        RECT  47.425 155.130 47.705 171.370 ;
        RECT  60.635 155.175 60.945 171.290 ;
        RECT  63.220 155.270 63.530 171.290 ;
        RECT  0.600 155.310 64.400 171.290 ;
        RECT  43.485 155.310 56.355 171.370 ;
        RECT  29.195 155.310 31.610 171.480 ;
        RECT  2.000 0.000 63.000 60.210 ;
        RECT  0.600 0.600 64.400 60.210 ;
        RECT  0.600 0.600 1.210 135.520 ;
        RECT  0.600 91.020 64.400 135.520 ;
        RECT  4.080 91.020 60.940 135.690 ;
        LAYER M3 ;
        RECT  0.600 247.660 25.790 248.740 ;
        RECT  0.600 247.660 25.470 249.400 ;
        RECT  28.830 247.660 64.400 248.740 ;
        RECT  29.150 247.660 29.470 249.400 ;
        RECT  31.880 247.660 64.400 249.400 ;
        RECT  0.600 124.090 64.400 129.850 ;
        RECT  4.040 123.970 60.900 135.790 ;
        RECT  1.640 124.090 63.600 135.790 ;
        RECT  1.810 124.090 2.830 154.520 ;
        RECT  1.640 155.040 63.600 171.560 ;
        RECT  1.640 183.580 63.600 185.950 ;
        RECT  2.790 155.040 63.600 200.820 ;
        RECT  4.860 124.090 63.600 200.820 ;
        RECT  1.640 196.170 63.600 200.820 ;
        RECT  0.600 0.600 64.400 60.480 ;
        RECT  2.000 0.000 63.000 88.700 ;
        RECT  0.600 0.600 1.480 91.220 ;
        RECT  0.600 90.750 64.400 91.220 ;
        LAYER TOP_M ;
        RECT  0.600 247.690 64.400 248.850 ;
        RECT  0.600 247.690 25.580 249.400 ;
        RECT  29.040 247.690 29.580 249.400 ;
        RECT  31.770 247.690 64.400 249.400 ;
        RECT  2.000 0.000 63.000 91.190 ;
        RECT  0.600 0.600 64.400 91.190 ;
    END
END pc3o02

MACRO pc3o01hv
    CLASS PAD ;
    FOREIGN pc3o01hv 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 65.000 BY 250.000 ;
    SYMMETRY X Y R90 ;
    SITE IOSite_c ;
    PIN PAD
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 55.440  LAYER TOP_M  ;
        ANTENNAPARTIALMETALSIDEAREA 287.938  LAYER M3  ;
        ANTENNAPARTIALMETALSIDEAREA 480.740  LAYER M2  ;
        ANTENNADIFFAREA 2657.280  LAYER TOP_M  ;
        ANTENNADIFFAREA 2657.280  LAYER M3  ;
        ANTENNADIFFAREA 1209.600  LAYER M2  ;
        ANTENNAPARTIALCUTAREA 632.318  LAYER TOP_V  ;
        ANTENNAPARTIALCUTAREA 349.898  LAYER V3  ;
        ANTENNAPARTIALCUTAREA 255.798  LAYER V2  ;
        PORT
        LAYER M3 ;
        RECT  26.310 249.580 28.310 250.000 ;
        LAYER M2 ;
        RECT  2.000 61.000 63.000 90.230 ;
        RECT  26.310 246.275 28.310 250.000 ;
        END
    END PAD
    PIN I
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 67.374  LAYER M1  ;
        ANTENNAPARTIALMETALSIDEAREA 81.652  LAYER M2  ;
        ANTENNAPARTIALMETALSIDEAREA 41.425  LAYER M3  ;
        ANTENNADIFFAREA 1.000  LAYER M3  ;
        ANTENNAPARTIALCUTAREA 0.203  LAYER V2  ;
        ANTENNAPARTIALCUTAREA 0.135  LAYER V3  ;
        ANTENNAGATEAREA 4.680  LAYER M2  ;
        ANTENNAGATEAREA 4.680  LAYER M3  ;
        PORT
        LAYER M3 ;
        RECT  30.310 249.580 31.040 250.000 ;
        LAYER M2 ;
        RECT  30.310 249.580 31.040 250.000 ;
        END
    END I
    PIN VDDO
        DIRECTION INOUT ;
        USE power ;
        PORT
        LAYER M3 ;
        RECT  64.200 192.330 65.000 200.640 ;
        RECT  0.000 201.660 65.000 221.520 ;
        RECT  0.000 222.720 65.000 246.820 ;
        RECT  0.000 192.330 0.800 200.640 ;
        LAYER M2 ;
        RECT  0.000 186.470 65.000 195.650 ;
        LAYER TOP_M ;
        RECT  0.000 195.170 65.000 200.640 ;
        RECT  0.000 201.660 65.000 221.520 ;
        RECT  0.000 222.720 65.000 246.820 ;
        END
    END VDDO
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        PORT
        LAYER M3 ;
        RECT  64.200 163.510 65.000 190.890 ;
        RECT  0.000 163.510 0.800 190.890 ;
        LAYER M2 ;
        RECT  0.000 172.080 65.000 183.060 ;
        LAYER TOP_M ;
        RECT  0.000 163.500 65.000 194.560 ;
        END
    END VDD
    PIN VSSO
        DIRECTION INOUT ;
        USE ground ;
        PORT
        LAYER M3 ;
        RECT  0.000 92.060 65.000 123.250 ;
        RECT  64.200 149.940 65.000 162.610 ;
        RECT  0.000 149.940 0.800 162.610 ;
        LAYER M2 ;
        RECT  0.000 147.040 65.000 154.520 ;
        LAYER TOP_M ;
        RECT  0.000 92.060 65.000 123.250 ;
        RECT  0.000 155.410 65.000 162.610 ;
        END
    END VSSO
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        PORT
        LAYER M3 ;
        RECT  64.200 130.690 65.000 148.880 ;
        RECT  0.000 130.690 0.800 148.880 ;
        LAYER M2 ;
        RECT  0.000 136.310 65.000 146.340 ;
        LAYER TOP_M ;
        RECT  0.000 123.850 65.000 154.560 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  2.000 0.000 63.000 250.000 ;
        RECT  0.000 88.990 65.000 130.360 ;
        RECT  0.000 136.510 65.000 157.550 ;
        RECT  0.300 158.930 64.700 159.230 ;
        RECT  0.300 159.530 64.700 159.830 ;
        RECT  0.300 160.130 64.700 160.430 ;
        RECT  0.300 160.730 64.700 161.030 ;
        RECT  0.300 161.330 64.700 161.630 ;
        RECT  0.300 161.910 64.700 162.190 ;
        RECT  0.300 162.490 64.700 162.770 ;
        RECT  0.300 163.070 64.700 163.350 ;
        RECT  0.300 163.650 64.700 163.950 ;
        RECT  0.300 164.250 64.700 164.550 ;
        RECT  0.300 164.850 64.700 165.150 ;
        RECT  0.300 165.450 64.700 165.750 ;
        RECT  0.300 166.050 64.700 166.350 ;
        RECT  0.300 166.650 64.700 166.960 ;
        RECT  0.300 167.260 64.700 167.560 ;
        RECT  0.300 167.860 64.700 168.160 ;
        RECT  0.000 169.150 65.000 197.240 ;
        RECT  0.600 0.600 64.400 250.000 ;
        RECT  0.000 198.470 65.000 250.000 ;
        LAYER M2 ;
        RECT  2.520 196.270 2.940 249.400 ;
        RECT  63.180 196.430 63.670 249.400 ;
        RECT  0.600 196.440 64.400 245.485 ;
        RECT  29.100 196.440 64.400 248.790 ;
        RECT  0.600 196.440 25.520 249.400 ;
        RECT  29.100 196.440 29.520 249.400 ;
        RECT  31.830 196.440 64.400 249.400 ;
        RECT  55.890 183.790 56.190 185.680 ;
        RECT  0.600 183.850 64.400 185.680 ;
        RECT  46.070 183.850 51.600 185.820 ;
        RECT  32.040 154.960 32.340 171.290 ;
        RECT  43.245 155.035 43.525 171.290 ;
        RECT  45.955 155.280 46.235 171.370 ;
        RECT  60.705 155.175 61.015 171.290 ;
        RECT  63.290 155.270 63.600 171.290 ;
        RECT  0.600 155.310 64.400 171.290 ;
        RECT  43.485 155.310 56.355 171.370 ;
        RECT  34.710 155.120 41.040 171.480 ;
        RECT  2.000 0.000 63.000 60.210 ;
        RECT  0.600 0.600 64.400 60.210 ;
        RECT  0.600 0.600 1.210 135.520 ;
        RECT  0.600 91.020 64.400 135.520 ;
        RECT  4.080 91.020 60.940 135.690 ;
        LAYER M3 ;
        RECT  0.600 247.660 25.790 248.740 ;
        RECT  0.600 247.660 25.470 249.400 ;
        RECT  28.830 247.660 64.400 248.740 ;
        RECT  29.150 247.660 29.470 249.400 ;
        RECT  31.880 247.660 64.400 249.400 ;
        RECT  4.040 123.870 60.900 200.820 ;
        RECT  0.600 124.090 64.400 129.850 ;
        RECT  1.640 124.090 63.600 135.790 ;
        RECT  1.810 124.090 2.830 154.520 ;
        RECT  1.640 155.040 63.600 171.560 ;
        RECT  1.640 183.580 63.600 185.950 ;
        RECT  2.520 155.040 63.600 200.820 ;
        RECT  4.040 124.090 63.600 200.820 ;
        RECT  1.640 196.170 63.600 200.820 ;
        RECT  0.600 0.600 64.400 60.480 ;
        RECT  2.000 0.000 63.000 88.700 ;
        RECT  0.600 0.600 1.480 91.220 ;
        RECT  0.600 90.750 64.400 91.220 ;
        LAYER TOP_M ;
        RECT  0.600 247.690 64.400 248.850 ;
        RECT  0.600 247.690 25.580 249.400 ;
        RECT  29.040 247.690 29.580 249.400 ;
        RECT  31.770 247.690 64.400 249.400 ;
        RECT  2.000 0.000 63.000 91.190 ;
        RECT  0.600 0.600 64.400 91.190 ;
    END
END pc3o01hv

MACRO pc3o01
    CLASS PAD ;
    FOREIGN pc3o01 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 65.000 BY 250.000 ;
    SYMMETRY X Y R90 ;
    SITE IOSite_c ;
    PIN PAD
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 55.440  LAYER TOP_M  ;
        ANTENNAPARTIALMETALSIDEAREA 287.938  LAYER M3  ;
        ANTENNAPARTIALMETALSIDEAREA 480.740  LAYER M2  ;
        ANTENNADIFFAREA 2657.280  LAYER TOP_M  ;
        ANTENNADIFFAREA 2657.280  LAYER M3  ;
        ANTENNADIFFAREA 1209.600  LAYER M2  ;
        ANTENNAPARTIALCUTAREA 632.318  LAYER TOP_V  ;
        ANTENNAPARTIALCUTAREA 349.898  LAYER V3  ;
        ANTENNAPARTIALCUTAREA 255.798  LAYER V2  ;
        PORT
        LAYER M3 ;
        RECT  26.310 249.580 28.310 250.000 ;
        LAYER M2 ;
        RECT  2.000 61.000 63.000 90.230 ;
        RECT  26.310 246.275 28.310 250.000 ;
        END
    END PAD
    PIN I
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 67.374  LAYER M1  ;
        ANTENNAPARTIALMETALSIDEAREA 81.652  LAYER M2  ;
        ANTENNAPARTIALMETALSIDEAREA 41.425  LAYER M3  ;
        ANTENNADIFFAREA 0.250  LAYER M3  ;
        ANTENNAPARTIALCUTAREA 0.270  LAYER V2  ;
        ANTENNAPARTIALCUTAREA 0.135  LAYER V3  ;
        ANTENNAGATEAREA 8.100  LAYER M2  ;
        ANTENNAGATEAREA 9.900  LAYER M3  ;
        PORT
        LAYER M3 ;
        RECT  30.310 249.580 31.040 250.000 ;
        LAYER M2 ;
        RECT  30.310 249.580 31.040 250.000 ;
        END
    END I
    PIN VDDO
        DIRECTION INOUT ;
        USE power ;
        PORT
        LAYER M3 ;
        RECT  64.200 192.330 65.000 200.640 ;
        RECT  0.000 201.660 65.000 221.520 ;
        RECT  0.000 222.720 65.000 246.820 ;
        RECT  0.000 192.330 0.800 200.640 ;
        LAYER M2 ;
        RECT  0.000 186.470 65.000 195.650 ;
        LAYER TOP_M ;
        RECT  0.000 195.170 65.000 200.640 ;
        RECT  0.000 201.660 65.000 221.520 ;
        RECT  0.000 222.720 65.000 246.820 ;
        END
    END VDDO
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        PORT
        LAYER M3 ;
        RECT  64.200 163.510 65.000 190.890 ;
        RECT  0.000 163.510 0.800 190.890 ;
        LAYER M2 ;
        RECT  0.000 172.080 65.000 183.060 ;
        LAYER TOP_M ;
        RECT  0.000 163.500 65.000 194.560 ;
        END
    END VDD
    PIN VSSO
        DIRECTION INOUT ;
        USE ground ;
        PORT
        LAYER M3 ;
        RECT  0.000 92.060 65.000 123.250 ;
        RECT  64.200 149.940 65.000 162.610 ;
        RECT  0.000 149.940 0.800 162.610 ;
        LAYER M2 ;
        RECT  0.000 147.040 65.000 154.520 ;
        LAYER TOP_M ;
        RECT  0.000 92.060 65.000 123.250 ;
        RECT  0.000 155.410 65.000 162.610 ;
        END
    END VSSO
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        PORT
        LAYER M3 ;
        RECT  64.200 130.690 65.000 148.880 ;
        RECT  0.000 130.690 0.800 148.880 ;
        LAYER M2 ;
        RECT  0.000 136.310 65.000 146.340 ;
        LAYER TOP_M ;
        RECT  0.000 123.850 65.000 154.560 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  2.000 0.000 63.000 250.000 ;
        RECT  0.000 88.990 65.000 130.360 ;
        RECT  0.000 136.510 65.000 157.550 ;
        RECT  0.300 158.930 64.700 159.230 ;
        RECT  0.300 159.530 64.700 159.830 ;
        RECT  0.300 160.130 64.700 160.430 ;
        RECT  0.300 160.730 64.700 161.030 ;
        RECT  0.300 161.330 64.700 161.630 ;
        RECT  0.300 161.910 64.700 162.190 ;
        RECT  0.300 162.490 64.700 162.770 ;
        RECT  0.300 163.070 64.700 163.350 ;
        RECT  0.300 163.650 64.700 163.950 ;
        RECT  0.300 164.250 64.700 164.550 ;
        RECT  0.300 164.850 64.700 165.150 ;
        RECT  0.300 165.450 64.700 165.750 ;
        RECT  0.300 166.050 64.700 166.350 ;
        RECT  0.300 166.650 64.700 166.960 ;
        RECT  0.300 167.260 64.700 167.560 ;
        RECT  0.300 167.860 64.700 168.160 ;
        RECT  0.000 169.150 65.000 197.240 ;
        RECT  0.600 0.600 64.400 250.000 ;
        RECT  0.000 198.470 65.000 250.000 ;
        LAYER M2 ;
        RECT  2.520 196.270 2.940 249.400 ;
        RECT  63.180 196.430 63.670 249.400 ;
        RECT  0.600 196.440 64.400 245.485 ;
        RECT  29.100 196.440 64.400 248.790 ;
        RECT  0.600 196.440 25.520 249.400 ;
        RECT  29.100 196.440 29.520 249.400 ;
        RECT  31.830 196.440 64.400 249.400 ;
        RECT  55.890 183.790 56.190 185.680 ;
        RECT  58.060 183.750 58.350 185.680 ;
        RECT  0.600 183.850 64.400 185.680 ;
        RECT  46.070 183.850 51.600 185.820 ;
        RECT  43.245 155.035 43.525 171.290 ;
        RECT  45.955 155.280 46.235 171.370 ;
        RECT  47.425 155.130 47.705 171.370 ;
        RECT  60.705 155.175 61.015 171.290 ;
        RECT  63.290 155.270 63.600 171.290 ;
        RECT  0.600 155.310 64.400 171.290 ;
        RECT  43.485 155.310 56.355 171.370 ;
        RECT  29.195 155.310 31.610 171.480 ;
        RECT  2.000 0.000 63.000 60.210 ;
        RECT  0.600 0.600 64.400 60.210 ;
        RECT  0.600 0.600 1.210 135.520 ;
        RECT  0.600 91.020 64.400 135.520 ;
        RECT  4.080 91.020 60.940 135.690 ;
        LAYER M3 ;
        RECT  0.600 247.660 25.790 248.740 ;
        RECT  0.600 247.660 25.470 249.400 ;
        RECT  28.830 247.660 64.400 248.740 ;
        RECT  29.150 247.660 29.470 249.400 ;
        RECT  31.880 247.660 64.400 249.400 ;
        RECT  4.040 123.870 60.900 200.820 ;
        RECT  0.600 124.090 64.400 129.850 ;
        RECT  1.640 124.090 63.600 135.790 ;
        RECT  1.810 124.090 2.830 154.520 ;
        RECT  1.640 155.040 63.600 171.560 ;
        RECT  1.640 183.580 63.600 185.950 ;
        RECT  2.520 155.040 63.600 200.820 ;
        RECT  4.040 124.090 63.600 200.820 ;
        RECT  1.640 196.170 63.600 200.820 ;
        RECT  0.600 0.600 64.400 60.480 ;
        RECT  2.000 0.000 63.000 88.700 ;
        RECT  0.600 0.600 1.480 91.220 ;
        RECT  0.600 90.750 64.400 91.220 ;
        LAYER TOP_M ;
        RECT  0.600 247.690 64.400 248.850 ;
        RECT  0.600 247.690 25.580 249.400 ;
        RECT  29.040 247.690 29.580 249.400 ;
        RECT  31.770 247.690 64.400 249.400 ;
        RECT  2.000 0.000 63.000 91.190 ;
        RECT  0.600 0.600 64.400 91.190 ;
    END
END pc3o01

MACRO pc3d31u
    CLASS PAD ;
    FOREIGN pc3d31u 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 65.000 BY 250.000 ;
    SYMMETRY X Y R90 ;
    SITE IOSite_c ;
    PIN PAD
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 55.440  LAYER TOP_M  ;
        ANTENNAPARTIALMETALSIDEAREA 287.938  LAYER M3  ;
        ANTENNAPARTIALMETALSIDEAREA 480.740  LAYER M2  ;
        ANTENNADIFFAREA 2657.280  LAYER TOP_M  ;
        ANTENNADIFFAREA 2657.280  LAYER M3  ;
        ANTENNADIFFAREA 1209.600  LAYER M2  ;
        ANTENNAPARTIALCUTAREA 632.318  LAYER TOP_V  ;
        ANTENNAPARTIALCUTAREA 349.898  LAYER V3  ;
        ANTENNAPARTIALCUTAREA 255.798  LAYER V2  ;
        PORT
        LAYER M3 ;
        RECT  24.870 249.580 26.870 250.000 ;
        LAYER M2 ;
        RECT  2.000 61.000 63.000 90.230 ;
        RECT  24.870 246.275 26.870 250.000 ;
        END
    END PAD
    PIN CIN
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 40.715  LAYER M3  ;
        ANTENNAPARTIALMETALSIDEAREA 104.781  LAYER M2  ;
        ANTENNAPARTIALMETALSIDEAREA 67.374  LAYER M1  ;
        ANTENNADIFFAREA 21.020  LAYER M3  ;
        ANTENNAPARTIALCUTAREA 0.203  LAYER V2  ;
        ANTENNAPARTIALCUTAREA 0.135  LAYER V3  ;
        PORT
        LAYER M3 ;
        RECT  28.870 249.580 29.600 250.000 ;
        LAYER M2 ;
        RECT  28.870 249.580 29.600 250.000 ;
        END
    END CIN
    PIN VDDO
        DIRECTION INOUT ;
        USE power ;
        PORT
        LAYER M3 ;
        RECT  64.200 192.330 65.000 200.640 ;
        RECT  0.000 201.660 65.000 221.520 ;
        RECT  0.000 222.720 65.000 246.820 ;
        RECT  0.000 192.330 0.800 200.640 ;
        LAYER M2 ;
        RECT  0.000 186.470 65.000 195.650 ;
        LAYER TOP_M ;
        RECT  0.000 195.170 65.000 200.640 ;
        RECT  0.000 201.660 65.000 221.520 ;
        RECT  0.000 222.720 65.000 246.820 ;
        END
    END VDDO
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        PORT
        LAYER M3 ;
        RECT  64.200 163.510 65.000 190.890 ;
        RECT  0.000 163.510 0.800 190.890 ;
        LAYER M2 ;
        RECT  0.000 172.080 65.000 183.060 ;
        LAYER TOP_M ;
        RECT  0.000 163.500 65.000 194.560 ;
        END
    END VDD
    PIN VSSO
        DIRECTION INOUT ;
        USE ground ;
        PORT
        LAYER M3 ;
        RECT  0.000 92.060 65.000 123.250 ;
        RECT  64.200 149.940 65.000 162.610 ;
        RECT  0.000 149.940 0.800 162.610 ;
        LAYER M2 ;
        RECT  0.000 147.040 65.000 154.520 ;
        LAYER TOP_M ;
        RECT  0.000 92.060 65.000 123.250 ;
        RECT  0.000 155.410 65.000 162.610 ;
        END
    END VSSO
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        PORT
        LAYER M3 ;
        RECT  64.200 130.690 65.000 148.880 ;
        RECT  0.000 130.690 0.800 148.880 ;
        LAYER M2 ;
        RECT  0.000 136.310 65.000 146.340 ;
        LAYER TOP_M ;
        RECT  0.000 123.850 65.000 154.560 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  2.000 0.000 63.000 250.000 ;
        RECT  0.000 88.990 65.000 130.360 ;
        RECT  0.000 136.510 65.000 157.550 ;
        RECT  0.315 158.150 64.700 158.460 ;
        RECT  0.300 158.930 64.700 159.230 ;
        RECT  0.300 159.530 64.700 159.830 ;
        RECT  0.300 160.130 64.700 160.430 ;
        RECT  0.300 160.730 64.700 161.030 ;
        RECT  0.300 161.330 64.700 161.630 ;
        RECT  0.300 161.910 64.700 162.190 ;
        RECT  0.300 162.490 64.700 162.770 ;
        RECT  0.300 163.070 64.700 163.350 ;
        RECT  0.300 163.650 64.700 163.950 ;
        RECT  0.300 164.250 64.700 164.550 ;
        RECT  0.300 164.850 64.700 165.150 ;
        RECT  0.300 165.450 64.700 165.750 ;
        RECT  0.300 166.050 64.700 166.350 ;
        RECT  0.300 166.650 64.700 166.960 ;
        RECT  0.300 167.260 64.700 167.560 ;
        RECT  0.300 167.860 64.700 168.160 ;
        RECT  0.000 169.150 65.000 197.240 ;
        RECT  0.600 0.600 64.400 250.000 ;
        RECT  0.000 198.470 65.000 250.000 ;
        LAYER M2 ;
        RECT  1.840 196.420 2.120 249.400 ;
        RECT  63.180 196.430 63.670 249.400 ;
        RECT  0.600 196.440 64.400 245.485 ;
        RECT  27.660 196.440 64.400 248.790 ;
        RECT  0.600 196.440 24.080 249.400 ;
        RECT  27.660 196.440 28.080 249.400 ;
        RECT  30.390 196.440 64.400 249.400 ;
        RECT  0.600 183.850 64.400 185.680 ;
        RECT  27.520 183.850 39.000 185.870 ;
        RECT  41.620 155.170 41.940 171.290 ;
        RECT  55.660 155.220 55.980 171.290 ;
        RECT  0.600 155.310 64.400 171.290 ;
        RECT  14.610 155.310 15.110 171.375 ;
        RECT  6.160 155.310 6.440 171.380 ;
        RECT  38.480 155.310 38.810 171.480 ;
        RECT  45.620 155.310 45.900 171.480 ;
        RECT  50.025 155.310 51.995 171.480 ;
        RECT  2.000 0.000 63.000 60.210 ;
        RECT  0.600 0.600 64.400 60.210 ;
        RECT  0.600 0.600 1.210 135.520 ;
        RECT  0.600 91.020 64.400 135.520 ;
        RECT  4.080 91.020 60.940 135.690 ;
        RECT  62.580 91.020 62.995 135.710 ;
        LAYER M3 ;
        RECT  0.600 247.660 24.350 248.740 ;
        RECT  0.600 247.660 24.030 249.400 ;
        RECT  27.390 247.660 64.400 248.740 ;
        RECT  27.710 247.660 28.030 249.400 ;
        RECT  30.440 247.660 64.400 249.400 ;
        RECT  0.600 124.090 64.400 129.850 ;
        RECT  1.640 124.090 63.600 135.790 ;
        RECT  1.810 124.090 2.830 154.520 ;
        RECT  4.040 123.970 60.900 171.560 ;
        RECT  1.640 155.040 63.600 171.560 ;
        RECT  1.640 183.580 63.600 185.950 ;
        RECT  5.490 124.090 63.600 200.820 ;
        RECT  1.640 196.170 63.600 200.820 ;
        RECT  56.930 123.970 57.210 201.060 ;
        RECT  0.600 0.600 64.400 60.480 ;
        RECT  2.000 0.000 63.000 88.700 ;
        RECT  0.600 0.600 1.480 91.220 ;
        RECT  0.600 90.750 64.400 91.220 ;
        LAYER TOP_M ;
        RECT  0.600 247.690 64.400 248.850 ;
        RECT  0.600 247.690 24.140 249.400 ;
        RECT  27.600 247.690 28.140 249.400 ;
        RECT  30.330 247.690 64.400 249.400 ;
        RECT  2.000 0.000 63.000 91.190 ;
        RECT  0.600 0.600 64.400 91.190 ;
    END
END pc3d31u

MACRO pc3d31d
    CLASS PAD ;
    FOREIGN pc3d31d 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 65.000 BY 250.000 ;
    SYMMETRY X Y R90 ;
    SITE IOSite_c ;
    PIN PAD
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 55.440  LAYER TOP_M  ;
        ANTENNAPARTIALMETALSIDEAREA 287.938  LAYER M3  ;
        ANTENNAPARTIALMETALSIDEAREA 480.740  LAYER M2  ;
        ANTENNADIFFAREA 2657.280  LAYER TOP_M  ;
        ANTENNADIFFAREA 2657.280  LAYER M3  ;
        ANTENNADIFFAREA 1209.600  LAYER M2  ;
        ANTENNAPARTIALCUTAREA 632.318  LAYER TOP_V  ;
        ANTENNAPARTIALCUTAREA 349.898  LAYER V3  ;
        ANTENNAPARTIALCUTAREA 255.798  LAYER V2  ;
        PORT
        LAYER M3 ;
        RECT  24.870 249.580 26.870 250.000 ;
        LAYER M2 ;
        RECT  2.000 61.000 63.000 90.230 ;
        RECT  24.870 246.275 26.870 250.000 ;
        END
    END PAD
    PIN CIN
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 40.715  LAYER M3  ;
        ANTENNAPARTIALMETALSIDEAREA 104.781  LAYER M2  ;
        ANTENNAPARTIALMETALSIDEAREA 67.374  LAYER M1  ;
        ANTENNADIFFAREA 21.020  LAYER M3  ;
        ANTENNAPARTIALCUTAREA 0.135  LAYER V3  ;
        ANTENNAPARTIALCUTAREA 0.203  LAYER V2  ;
        PORT
        LAYER M3 ;
        RECT  28.870 249.580 29.600 250.000 ;
        LAYER M2 ;
        RECT  28.870 249.580 29.600 250.000 ;
        END
    END CIN
    PIN VDDO
        DIRECTION INOUT ;
        USE power ;
        PORT
        LAYER M3 ;
        RECT  64.200 192.330 65.000 200.640 ;
        RECT  0.000 201.660 65.000 221.520 ;
        RECT  0.000 222.720 65.000 246.820 ;
        RECT  0.000 192.330 0.800 200.640 ;
        LAYER M2 ;
        RECT  0.000 186.470 65.000 195.650 ;
        LAYER TOP_M ;
        RECT  0.000 195.170 65.000 200.640 ;
        RECT  0.000 201.660 65.000 221.520 ;
        RECT  0.000 222.720 65.000 246.820 ;
        END
    END VDDO
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        PORT
        LAYER M3 ;
        RECT  64.200 163.510 65.000 190.890 ;
        RECT  0.000 163.510 0.800 190.890 ;
        LAYER M2 ;
        RECT  0.000 172.080 65.000 183.060 ;
        LAYER TOP_M ;
        RECT  0.000 163.500 65.000 194.560 ;
        END
    END VDD
    PIN VSSO
        DIRECTION INOUT ;
        USE ground ;
        PORT
        LAYER M3 ;
        RECT  0.000 92.060 65.000 123.250 ;
        RECT  64.200 149.940 65.000 162.610 ;
        RECT  0.000 149.940 0.800 162.610 ;
        LAYER M2 ;
        RECT  0.000 147.040 65.000 154.520 ;
        LAYER TOP_M ;
        RECT  0.000 92.060 65.000 123.250 ;
        RECT  0.000 155.410 65.000 162.610 ;
        END
    END VSSO
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        PORT
        LAYER M3 ;
        RECT  64.200 130.690 65.000 148.880 ;
        RECT  0.000 130.690 0.800 148.880 ;
        LAYER M2 ;
        RECT  0.000 136.310 65.000 146.340 ;
        LAYER TOP_M ;
        RECT  0.000 123.850 65.000 154.560 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  2.000 0.000 63.000 250.000 ;
        RECT  0.000 88.990 65.000 130.360 ;
        RECT  0.000 136.510 65.000 157.550 ;
        RECT  0.315 158.150 64.700 158.460 ;
        RECT  0.300 158.930 64.700 159.230 ;
        RECT  0.300 159.530 64.700 159.830 ;
        RECT  0.300 160.130 64.700 160.430 ;
        RECT  0.300 160.730 64.700 161.030 ;
        RECT  0.300 161.330 64.700 161.630 ;
        RECT  0.300 161.910 64.700 162.190 ;
        RECT  0.300 162.490 64.700 162.770 ;
        RECT  0.300 163.070 64.700 163.350 ;
        RECT  0.300 163.650 64.700 163.950 ;
        RECT  0.300 164.250 64.700 164.550 ;
        RECT  0.300 164.850 64.700 165.150 ;
        RECT  0.300 165.450 64.700 165.750 ;
        RECT  0.300 166.050 64.700 166.350 ;
        RECT  0.300 166.650 64.700 166.960 ;
        RECT  0.300 167.260 64.700 167.560 ;
        RECT  0.300 167.860 64.700 168.160 ;
        RECT  0.000 169.150 65.000 197.240 ;
        RECT  0.600 0.600 64.400 250.000 ;
        RECT  0.000 198.470 65.000 250.000 ;
        LAYER M2 ;
        RECT  1.840 196.420 2.120 249.400 ;
        RECT  63.180 196.430 63.670 249.400 ;
        RECT  0.600 196.440 64.400 245.485 ;
        RECT  27.660 196.440 64.400 248.790 ;
        RECT  0.600 196.440 24.080 249.400 ;
        RECT  27.660 196.440 28.080 249.400 ;
        RECT  30.390 196.440 64.400 249.400 ;
        RECT  0.600 183.850 64.400 185.680 ;
        RECT  27.520 183.850 39.000 185.870 ;
        RECT  41.620 155.170 41.940 171.290 ;
        RECT  48.725 155.130 50.965 171.290 ;
        RECT  51.905 155.300 52.215 171.290 ;
        RECT  55.660 155.220 55.980 171.290 ;
        RECT  0.600 155.310 64.400 171.290 ;
        RECT  6.160 155.310 6.440 171.380 ;
        RECT  38.480 155.310 38.810 171.480 ;
        RECT  45.620 155.310 45.900 171.480 ;
        RECT  50.025 155.310 51.995 171.480 ;
        RECT  2.000 0.000 63.000 60.210 ;
        RECT  0.600 0.600 64.400 60.210 ;
        RECT  0.600 0.600 1.210 135.520 ;
        RECT  0.600 91.020 64.400 135.520 ;
        RECT  4.080 91.020 60.940 135.690 ;
        RECT  62.580 91.020 62.995 135.710 ;
        LAYER M3 ;
        RECT  0.600 247.660 24.350 248.740 ;
        RECT  0.600 247.660 24.030 249.400 ;
        RECT  27.390 247.660 64.400 248.740 ;
        RECT  27.710 247.660 28.030 249.400 ;
        RECT  30.440 247.660 64.400 249.400 ;
        RECT  0.600 124.090 64.400 129.850 ;
        RECT  1.640 124.090 63.600 135.790 ;
        RECT  1.810 124.090 2.830 154.520 ;
        RECT  4.040 123.970 60.900 171.560 ;
        RECT  1.640 155.040 63.600 171.560 ;
        RECT  1.640 183.580 63.600 185.950 ;
        RECT  5.490 124.090 63.600 200.820 ;
        RECT  1.640 196.170 63.600 200.820 ;
        RECT  56.930 123.970 57.210 201.060 ;
        RECT  0.600 0.600 64.400 60.480 ;
        RECT  2.000 0.000 63.000 88.700 ;
        RECT  0.600 0.600 1.480 91.220 ;
        RECT  0.600 90.750 64.400 91.220 ;
        LAYER TOP_M ;
        RECT  0.600 247.690 64.400 248.850 ;
        RECT  0.600 247.690 24.140 249.400 ;
        RECT  27.600 247.690 28.140 249.400 ;
        RECT  30.330 247.690 64.400 249.400 ;
        RECT  2.000 0.000 63.000 91.190 ;
        RECT  0.600 0.600 64.400 91.190 ;
    END
END pc3d31d

MACRO pc3d31
    CLASS PAD ;
    FOREIGN pc3d31 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 65.000 BY 250.000 ;
    SYMMETRY X Y R90 ;
    SITE IOSite_c ;
    PIN PAD
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 55.440  LAYER TOP_M  ;
        ANTENNAPARTIALMETALSIDEAREA 287.938  LAYER M3  ;
        ANTENNAPARTIALMETALSIDEAREA 480.740  LAYER M2  ;
        ANTENNADIFFAREA 2657.280  LAYER TOP_M  ;
        ANTENNADIFFAREA 2657.280  LAYER M3  ;
        ANTENNADIFFAREA 1209.600  LAYER M2  ;
        ANTENNAPARTIALCUTAREA 632.318  LAYER TOP_V  ;
        ANTENNAPARTIALCUTAREA 349.898  LAYER V3  ;
        ANTENNAPARTIALCUTAREA 255.798  LAYER V2  ;
        PORT
        LAYER M3 ;
        RECT  24.870 249.580 26.870 250.000 ;
        LAYER M2 ;
        RECT  2.000 61.000 63.000 90.230 ;
        RECT  24.870 246.275 26.870 250.000 ;
        END
    END PAD
    PIN CIN
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 40.715  LAYER M3  ;
        ANTENNAPARTIALMETALSIDEAREA 104.781  LAYER M2  ;
        ANTENNAPARTIALMETALSIDEAREA 67.374  LAYER M1  ;
        ANTENNADIFFAREA 21.020  LAYER M3  ;
        ANTENNAPARTIALCUTAREA 0.203  LAYER V2  ;
        ANTENNAPARTIALCUTAREA 0.135  LAYER V3  ;
        PORT
        LAYER M3 ;
        RECT  28.870 249.580 29.600 250.000 ;
        LAYER M2 ;
        RECT  28.870 249.580 29.600 250.000 ;
        END
    END CIN
    PIN VDDO
        DIRECTION INOUT ;
        USE power ;
        PORT
        LAYER M3 ;
        RECT  64.200 192.330 65.000 200.640 ;
        RECT  0.000 201.660 65.000 221.520 ;
        RECT  0.000 222.720 65.000 246.820 ;
        RECT  0.000 192.330 0.800 200.640 ;
        LAYER M2 ;
        RECT  0.000 186.470 65.000 195.650 ;
        LAYER TOP_M ;
        RECT  0.000 195.170 65.000 200.640 ;
        RECT  0.000 201.660 65.000 221.520 ;
        RECT  0.000 222.720 65.000 246.820 ;
        END
    END VDDO
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        PORT
        LAYER M3 ;
        RECT  64.200 163.510 65.000 190.890 ;
        RECT  0.000 163.510 0.800 190.890 ;
        LAYER M2 ;
        RECT  0.000 172.080 65.000 183.060 ;
        LAYER TOP_M ;
        RECT  0.000 163.500 65.000 194.560 ;
        END
    END VDD
    PIN VSSO
        DIRECTION INOUT ;
        USE ground ;
        PORT
        LAYER M3 ;
        RECT  0.000 92.060 65.000 123.250 ;
        RECT  64.200 149.940 65.000 162.610 ;
        RECT  0.000 149.940 0.800 162.610 ;
        LAYER M2 ;
        RECT  0.000 147.040 65.000 154.520 ;
        LAYER TOP_M ;
        RECT  0.000 92.060 65.000 123.250 ;
        RECT  0.000 155.410 65.000 162.610 ;
        END
    END VSSO
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        PORT
        LAYER M3 ;
        RECT  64.200 130.690 65.000 148.880 ;
        RECT  0.000 130.690 0.800 148.880 ;
        LAYER M2 ;
        RECT  0.000 136.310 65.000 146.340 ;
        LAYER TOP_M ;
        RECT  0.000 123.850 65.000 154.560 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  2.000 0.000 63.000 250.000 ;
        RECT  0.000 88.990 65.000 130.360 ;
        RECT  0.000 136.510 65.000 157.550 ;
        RECT  0.315 158.150 64.700 158.460 ;
        RECT  0.300 158.930 64.700 159.230 ;
        RECT  0.300 159.530 64.700 159.830 ;
        RECT  0.300 160.130 64.700 160.430 ;
        RECT  0.300 160.730 64.700 161.030 ;
        RECT  0.300 161.330 64.700 161.630 ;
        RECT  0.300 161.910 64.700 162.190 ;
        RECT  0.300 162.490 64.700 162.770 ;
        RECT  0.300 163.070 64.700 163.350 ;
        RECT  0.300 163.650 64.700 163.950 ;
        RECT  0.300 164.250 64.700 164.550 ;
        RECT  0.300 164.850 64.700 165.150 ;
        RECT  0.300 165.450 64.700 165.750 ;
        RECT  0.300 166.050 64.700 166.350 ;
        RECT  0.300 166.650 64.700 166.960 ;
        RECT  0.300 167.260 64.700 167.560 ;
        RECT  0.300 167.860 64.700 168.160 ;
        RECT  0.000 169.150 65.000 197.240 ;
        RECT  0.600 0.600 64.400 250.000 ;
        RECT  0.000 198.470 65.000 250.000 ;
        LAYER M2 ;
        RECT  1.840 196.420 2.120 249.400 ;
        RECT  63.180 196.430 63.670 249.400 ;
        RECT  0.600 196.440 64.400 245.485 ;
        RECT  27.660 196.440 64.400 248.790 ;
        RECT  0.600 196.440 24.080 249.400 ;
        RECT  27.660 196.440 28.080 249.400 ;
        RECT  30.390 196.440 64.400 249.400 ;
        RECT  0.600 183.850 64.400 185.680 ;
        RECT  27.520 183.850 39.000 185.870 ;
        RECT  41.620 155.170 41.940 171.290 ;
        RECT  55.660 155.220 55.980 171.290 ;
        RECT  0.600 155.310 64.400 171.290 ;
        RECT  6.160 155.310 6.440 171.380 ;
        RECT  38.480 155.310 38.810 171.480 ;
        RECT  45.620 155.310 45.900 171.480 ;
        RECT  50.025 155.310 51.995 171.480 ;
        RECT  2.000 0.000 63.000 60.210 ;
        RECT  0.600 0.600 64.400 60.210 ;
        RECT  0.600 0.600 1.210 135.520 ;
        RECT  0.600 91.020 64.400 135.520 ;
        RECT  4.080 91.020 60.940 135.690 ;
        RECT  62.580 91.020 62.995 135.710 ;
        LAYER M3 ;
        RECT  0.600 247.660 24.350 248.740 ;
        RECT  0.600 247.660 24.030 249.400 ;
        RECT  27.390 247.660 64.400 248.740 ;
        RECT  27.710 247.660 28.030 249.400 ;
        RECT  30.440 247.660 64.400 249.400 ;
        RECT  0.600 124.090 64.400 129.850 ;
        RECT  1.640 124.090 63.600 135.790 ;
        RECT  1.810 124.090 2.830 154.520 ;
        RECT  4.040 123.970 60.900 171.560 ;
        RECT  1.640 155.040 63.600 171.560 ;
        RECT  1.640 183.580 63.600 185.950 ;
        RECT  5.490 124.090 63.600 200.820 ;
        RECT  1.640 196.170 63.600 200.820 ;
        RECT  56.930 123.970 57.210 201.060 ;
        RECT  0.600 0.600 64.400 60.480 ;
        RECT  2.000 0.000 63.000 88.700 ;
        RECT  0.600 0.600 1.480 91.220 ;
        RECT  0.600 90.750 64.400 91.220 ;
        LAYER TOP_M ;
        RECT  0.600 247.690 64.400 248.850 ;
        RECT  0.600 247.690 24.140 249.400 ;
        RECT  27.600 247.690 28.140 249.400 ;
        RECT  30.330 247.690 64.400 249.400 ;
        RECT  2.000 0.000 63.000 91.190 ;
        RECT  0.600 0.600 64.400 91.190 ;
    END
END pc3d31

MACRO pc3d21u
    CLASS PAD ;
    FOREIGN pc3d21u 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 65.000 BY 250.000 ;
    SYMMETRY X Y R90 ;
    SITE IOSite_c ;
    PIN PAD
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 55.440  LAYER TOP_M  ;
        ANTENNAPARTIALMETALSIDEAREA 287.938  LAYER M3  ;
        ANTENNAPARTIALMETALSIDEAREA 480.740  LAYER M2  ;
        ANTENNADIFFAREA 2657.280  LAYER TOP_M  ;
        ANTENNADIFFAREA 2657.280  LAYER M3  ;
        ANTENNADIFFAREA 1209.600  LAYER M2  ;
        ANTENNAPARTIALCUTAREA 255.798  LAYER V2  ;
        ANTENNAPARTIALCUTAREA 632.318  LAYER TOP_V  ;
        ANTENNAPARTIALCUTAREA 349.898  LAYER V3  ;
        PORT
        LAYER M2 ;
        RECT  2.000 61.000 63.000 90.230 ;
        RECT  24.870 246.275 26.870 250.000 ;
        LAYER M3 ;
        RECT  24.870 249.580 26.870 250.000 ;
        END
    END PAD
    PIN CIN
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 67.374  LAYER M1  ;
        ANTENNAPARTIALMETALSIDEAREA 188.733  LAYER M2  ;
        ANTENNAPARTIALMETALSIDEAREA 40.715  LAYER M3  ;
        ANTENNADIFFAREA 21.020  LAYER M3  ;
        ANTENNADIFFAREA 21.020  LAYER M2  ;
        ANTENNAPARTIALCUTAREA 0.270  LAYER V2  ;
        ANTENNAPARTIALCUTAREA 0.203  LAYER V3  ;
        PORT
        LAYER M2 ;
        RECT  28.870 249.580 29.600 250.000 ;
        LAYER M3 ;
        RECT  28.870 249.580 29.600 250.000 ;
        END
    END CIN
    PIN VDDO
        DIRECTION INOUT ;
        USE power ;
        PORT
        LAYER TOP_M ;
        RECT  0.000 195.170 65.000 200.640 ;
        RECT  0.000 201.660 65.000 221.520 ;
        RECT  0.000 222.720 65.000 246.820 ;
        LAYER M2 ;
        RECT  0.000 186.470 65.000 195.650 ;
        LAYER M3 ;
        RECT  64.200 192.330 65.000 200.640 ;
        RECT  0.000 201.660 65.000 221.520 ;
        RECT  0.000 222.720 65.000 246.820 ;
        RECT  0.000 192.330 0.800 200.640 ;
        END
    END VDDO
    PIN VSSO
        DIRECTION INOUT ;
        USE ground ;
        PORT
        LAYER TOP_M ;
        RECT  0.000 92.060 65.000 123.250 ;
        RECT  0.000 155.410 65.000 162.610 ;
        LAYER M2 ;
        RECT  0.000 147.040 65.000 154.520 ;
        LAYER M3 ;
        RECT  0.000 92.060 65.000 123.250 ;
        RECT  64.200 149.940 65.000 162.610 ;
        RECT  0.000 149.940 0.800 162.610 ;
        END
    END VSSO
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        PORT
        LAYER TOP_M ;
        RECT  0.000 123.850 65.000 154.560 ;
        LAYER M2 ;
        RECT  0.000 136.310 65.000 146.340 ;
        LAYER M3 ;
        RECT  64.200 130.690 65.000 148.880 ;
        RECT  0.000 130.690 0.800 148.880 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        PORT
        LAYER TOP_M ;
        RECT  0.000 163.500 65.000 194.560 ;
        LAYER M2 ;
        RECT  0.000 172.080 65.000 183.060 ;
        LAYER M3 ;
        RECT  64.200 163.510 65.000 190.890 ;
        RECT  0.000 163.510 0.800 190.890 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.000 0.000 63.000 250.000 ;
        RECT  0.000 88.990 65.000 130.360 ;
        RECT  0.000 136.510 65.000 157.550 ;
        RECT  0.315 158.150 64.700 158.460 ;
        RECT  0.300 158.930 64.700 159.230 ;
        RECT  0.300 159.530 64.700 159.830 ;
        RECT  0.300 160.130 64.700 160.430 ;
        RECT  0.300 160.730 64.700 161.030 ;
        RECT  0.300 161.330 64.700 161.630 ;
        RECT  0.300 161.910 64.700 162.190 ;
        RECT  0.300 162.490 64.700 162.770 ;
        RECT  0.300 163.070 64.700 163.350 ;
        RECT  0.300 163.650 64.700 163.950 ;
        RECT  0.300 164.250 64.700 164.550 ;
        RECT  0.300 164.850 64.700 165.150 ;
        RECT  0.300 165.450 64.700 165.750 ;
        RECT  0.300 166.050 64.700 166.350 ;
        RECT  0.300 166.650 64.700 166.960 ;
        RECT  0.300 167.260 64.700 167.560 ;
        RECT  0.300 167.860 64.700 168.160 ;
        RECT  0.000 169.150 65.000 197.240 ;
        RECT  0.600 0.600 64.400 250.000 ;
        RECT  0.000 198.470 65.000 250.000 ;
        LAYER M2 ;
        RECT  1.840 196.420 2.120 249.400 ;
        RECT  63.180 196.430 63.670 249.400 ;
        RECT  0.600 196.440 64.400 245.485 ;
        RECT  27.660 196.440 64.400 248.790 ;
        RECT  0.600 196.440 24.080 249.400 ;
        RECT  27.660 196.440 28.080 249.400 ;
        RECT  30.390 196.440 64.400 249.400 ;
        RECT  0.600 183.850 64.400 185.680 ;
        RECT  32.400 155.220 32.720 171.290 ;
        RECT  0.600 155.310 64.400 171.290 ;
        RECT  13.770 155.310 14.270 171.375 ;
        RECT  6.160 155.310 6.440 171.380 ;
        RECT  45.210 155.310 45.490 171.480 ;
        RECT  50.025 155.310 51.995 171.480 ;
        RECT  2.000 0.000 63.000 60.210 ;
        RECT  0.600 0.600 64.400 60.210 ;
        RECT  0.600 0.600 1.210 135.520 ;
        RECT  0.600 91.020 64.400 135.520 ;
        RECT  4.080 91.020 60.940 135.690 ;
        RECT  62.580 91.020 62.995 135.710 ;
        LAYER M3 ;
        RECT  0.600 247.660 24.350 248.740 ;
        RECT  0.600 247.660 24.030 249.400 ;
        RECT  27.390 247.660 64.400 248.740 ;
        RECT  27.710 247.660 28.030 249.400 ;
        RECT  30.440 247.660 64.400 249.400 ;
        RECT  0.600 124.090 64.400 129.850 ;
        RECT  1.640 124.090 63.600 135.790 ;
        RECT  1.810 124.090 2.830 154.520 ;
        RECT  4.040 123.970 60.900 171.560 ;
        RECT  1.640 155.040 63.600 171.560 ;
        RECT  1.640 183.580 63.600 185.950 ;
        RECT  5.490 124.090 63.600 200.820 ;
        RECT  1.640 196.170 63.600 200.820 ;
        RECT  56.930 123.970 57.210 201.060 ;
        RECT  0.600 0.600 64.400 60.480 ;
        RECT  2.000 0.000 63.000 88.700 ;
        RECT  0.600 0.600 1.480 91.220 ;
        RECT  0.600 90.750 64.400 91.220 ;
        LAYER TOP_M ;
        RECT  0.600 247.690 64.400 248.850 ;
        RECT  0.600 247.690 24.140 249.400 ;
        RECT  27.600 247.690 28.140 249.400 ;
        RECT  30.330 247.690 64.400 249.400 ;
        RECT  2.000 0.000 63.000 91.190 ;
        RECT  0.600 0.600 64.400 91.190 ;
    END
END pc3d21u

MACRO pc3d21eu
    CLASS PAD ;
    FOREIGN pc3d21eu 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 65.000 BY 250.000 ;
    SYMMETRY X Y R90 ;
    SITE IOSite_c ;
    PIN RENB
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 67.310  LAYER M1  ;
        ANTENNAPARTIALMETALSIDEAREA 80.528  LAYER M2  ;
        ANTENNAPARTIALMETALSIDEAREA 40.105  LAYER M3  ;
        ANTENNADIFFAREA 1.000  LAYER M3  ;
        ANTENNAPARTIALCUTAREA 0.135  LAYER V3  ;
        ANTENNAPARTIALCUTAREA 0.203  LAYER V2  ;
        ANTENNAGATEAREA 5.760  LAYER M2  ;
        ANTENNAGATEAREA 6.316  LAYER M3  ;
        PORT
        LAYER M2 ;
        RECT  29.900 249.620 30.630 250.000 ;
        LAYER M3 ;
        RECT  29.900 249.620 30.630 250.000 ;
        END
    END RENB
    PIN PAD
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 55.440  LAYER TOP_M  ;
        ANTENNAPARTIALMETALSIDEAREA 287.938  LAYER M3  ;
        ANTENNAPARTIALMETALSIDEAREA 480.740  LAYER M2  ;
        ANTENNADIFFAREA 2657.280  LAYER TOP_M  ;
        ANTENNADIFFAREA 2657.280  LAYER M3  ;
        ANTENNADIFFAREA 1209.600  LAYER M2  ;
        ANTENNAPARTIALCUTAREA 255.798  LAYER V2  ;
        ANTENNAPARTIALCUTAREA 632.318  LAYER TOP_V  ;
        ANTENNAPARTIALCUTAREA 349.898  LAYER V3  ;
        PORT
        LAYER M2 ;
        RECT  2.000 61.000 63.000 90.230 ;
        RECT  24.870 246.275 26.870 250.000 ;
        LAYER M3 ;
        RECT  24.870 249.580 26.870 250.000 ;
        END
    END PAD
    PIN CIN
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 67.374  LAYER M1  ;
        ANTENNAPARTIALMETALSIDEAREA 184.673  LAYER M2  ;
        ANTENNAPARTIALMETALSIDEAREA 40.715  LAYER M3  ;
        ANTENNADIFFAREA 21.020  LAYER M2  ;
        ANTENNADIFFAREA 21.020  LAYER M3  ;
        ANTENNAPARTIALCUTAREA 0.270  LAYER V2  ;
        ANTENNAPARTIALCUTAREA 0.203  LAYER V3  ;
        PORT
        LAYER M2 ;
        RECT  28.870 249.620 29.600 250.000 ;
        LAYER M3 ;
        RECT  28.870 249.620 29.600 250.000 ;
        END
    END CIN
    PIN VDDO
        DIRECTION INOUT ;
        USE power ;
        PORT
        LAYER TOP_M ;
        RECT  0.000 195.170 65.000 200.640 ;
        RECT  0.000 201.660 65.000 221.520 ;
        RECT  0.000 222.720 65.000 246.820 ;
        LAYER M2 ;
        RECT  0.000 186.470 65.000 195.650 ;
        LAYER M3 ;
        RECT  64.200 192.330 65.000 200.640 ;
        RECT  0.000 201.660 65.000 221.520 ;
        RECT  0.000 222.720 65.000 246.820 ;
        RECT  0.000 192.330 0.800 200.640 ;
        END
    END VDDO
    PIN VSSO
        DIRECTION INOUT ;
        USE ground ;
        PORT
        LAYER TOP_M ;
        RECT  0.000 92.060 65.000 123.250 ;
        RECT  0.000 155.410 65.000 162.610 ;
        LAYER M2 ;
        RECT  0.000 147.040 65.000 154.520 ;
        LAYER M3 ;
        RECT  0.000 92.060 65.000 123.250 ;
        RECT  64.200 149.940 65.000 162.610 ;
        RECT  0.000 149.940 0.800 162.610 ;
        END
    END VSSO
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        PORT
        LAYER TOP_M ;
        RECT  0.000 123.850 65.000 154.560 ;
        LAYER M2 ;
        RECT  0.000 136.310 65.000 146.340 ;
        LAYER M3 ;
        RECT  64.200 130.690 65.000 148.880 ;
        RECT  0.000 130.690 0.800 148.880 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        PORT
        LAYER TOP_M ;
        RECT  0.000 163.500 65.000 194.560 ;
        LAYER M2 ;
        RECT  0.000 172.080 65.000 183.060 ;
        LAYER M3 ;
        RECT  64.200 163.510 65.000 190.890 ;
        RECT  0.000 163.510 0.800 190.890 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.000 0.000 63.000 250.000 ;
        RECT  0.000 88.990 65.000 130.360 ;
        RECT  0.000 136.510 65.000 157.550 ;
        RECT  0.300 158.930 64.700 159.230 ;
        RECT  0.300 159.530 64.700 159.830 ;
        RECT  0.300 160.130 64.700 160.430 ;
        RECT  0.300 160.730 64.700 161.030 ;
        RECT  0.300 161.330 64.700 161.630 ;
        RECT  0.300 161.910 64.700 162.190 ;
        RECT  0.300 162.490 64.700 162.770 ;
        RECT  0.300 163.070 64.700 163.350 ;
        RECT  0.300 163.650 64.700 163.950 ;
        RECT  0.300 164.250 64.700 164.550 ;
        RECT  0.300 164.850 64.700 165.150 ;
        RECT  0.300 165.450 64.700 165.750 ;
        RECT  0.300 166.050 64.700 166.350 ;
        RECT  0.300 166.650 64.700 166.960 ;
        RECT  0.300 167.260 64.700 167.560 ;
        RECT  0.300 167.860 64.700 168.160 ;
        RECT  0.000 169.150 65.000 197.240 ;
        RECT  0.600 0.600 64.400 250.000 ;
        RECT  0.000 198.470 65.000 250.000 ;
        LAYER M2 ;
        RECT  1.840 196.420 2.120 249.400 ;
        RECT  63.180 196.430 63.670 249.400 ;
        RECT  0.600 196.440 64.400 245.485 ;
        RECT  27.660 196.440 64.400 248.830 ;
        RECT  0.600 196.440 24.080 249.400 ;
        RECT  27.660 196.440 28.080 249.400 ;
        RECT  31.420 196.440 64.400 249.400 ;
        RECT  57.720 183.660 58.680 185.870 ;
        RECT  0.600 183.850 64.400 185.680 ;
        RECT  57.500 183.850 58.880 185.870 ;
        RECT  32.400 155.220 32.720 171.290 ;
        RECT  0.600 155.310 64.400 171.290 ;
        RECT  6.160 155.310 6.440 171.380 ;
        RECT  38.250 155.310 40.585 171.460 ;
        RECT  41.815 155.310 42.200 171.480 ;
        RECT  45.210 155.310 45.490 171.480 ;
        RECT  50.025 155.310 51.995 171.480 ;
        RECT  2.000 0.000 63.000 60.210 ;
        RECT  0.600 0.600 64.400 60.210 ;
        RECT  0.600 0.600 1.210 135.520 ;
        RECT  0.600 91.020 64.400 135.520 ;
        RECT  4.080 91.020 60.940 135.690 ;
        RECT  62.580 91.020 62.995 135.710 ;
        LAYER M3 ;
        RECT  0.600 247.660 24.350 248.740 ;
        RECT  0.600 247.660 24.030 249.400 ;
        RECT  27.390 247.660 64.400 248.740 ;
        RECT  27.710 247.660 64.400 248.780 ;
        RECT  27.710 247.660 28.030 249.400 ;
        RECT  31.470 247.660 64.400 249.400 ;
        RECT  0.600 124.090 64.400 129.850 ;
        RECT  1.640 124.090 63.600 135.790 ;
        RECT  1.810 124.090 2.830 154.520 ;
        RECT  4.040 123.970 60.900 171.560 ;
        RECT  1.640 155.040 63.600 171.560 ;
        RECT  1.640 183.580 63.600 185.950 ;
        RECT  5.490 124.090 63.600 200.820 ;
        RECT  1.640 196.170 63.600 200.820 ;
        RECT  56.930 123.970 57.210 201.060 ;
        RECT  57.815 123.970 58.100 201.060 ;
        RECT  0.600 0.600 64.400 60.480 ;
        RECT  2.000 0.000 63.000 88.700 ;
        RECT  0.600 0.600 1.480 91.220 ;
        RECT  0.600 90.750 64.400 91.220 ;
        LAYER TOP_M ;
        RECT  0.600 247.690 64.400 248.850 ;
        RECT  27.600 247.690 64.400 248.890 ;
        RECT  0.600 247.690 24.140 249.400 ;
        RECT  27.600 247.690 28.140 249.400 ;
        RECT  31.360 247.690 64.400 249.400 ;
        RECT  2.000 0.000 63.000 91.190 ;
        RECT  0.600 0.600 64.400 91.190 ;
    END
END pc3d21eu

MACRO pc3d21d
    CLASS PAD ;
    FOREIGN pc3d21d 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 65.000 BY 250.000 ;
    SYMMETRY X Y R90 ;
    SITE IOSite_c ;
    PIN PAD
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 55.440  LAYER TOP_M  ;
        ANTENNAPARTIALMETALSIDEAREA 287.938  LAYER M3  ;
        ANTENNAPARTIALMETALSIDEAREA 480.740  LAYER M2  ;
        ANTENNADIFFAREA 2657.280  LAYER TOP_M  ;
        ANTENNADIFFAREA 2657.280  LAYER M3  ;
        ANTENNADIFFAREA 1209.600  LAYER M2  ;
        ANTENNAPARTIALCUTAREA 255.798  LAYER V2  ;
        ANTENNAPARTIALCUTAREA 632.318  LAYER TOP_V  ;
        ANTENNAPARTIALCUTAREA 349.898  LAYER V3  ;
        PORT
        LAYER M2 ;
        RECT  2.000 61.000 63.000 90.230 ;
        RECT  24.870 246.275 26.870 250.000 ;
        LAYER M3 ;
        RECT  24.870 249.580 26.870 250.000 ;
        END
    END PAD
    PIN CIN
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 67.374  LAYER M1  ;
        ANTENNAPARTIALMETALSIDEAREA 188.733  LAYER M2  ;
        ANTENNAPARTIALMETALSIDEAREA 40.715  LAYER M3  ;
        ANTENNADIFFAREA 21.020  LAYER M3  ;
        ANTENNADIFFAREA 21.020  LAYER M2  ;
        ANTENNAPARTIALCUTAREA 0.270  LAYER V2  ;
        ANTENNAPARTIALCUTAREA 0.203  LAYER V3  ;
        PORT
        LAYER M2 ;
        RECT  28.870 249.580 29.600 250.000 ;
        LAYER M3 ;
        RECT  28.870 249.580 29.600 250.000 ;
        END
    END CIN
    PIN VDDO
        DIRECTION INOUT ;
        USE power ;
        PORT
        LAYER TOP_M ;
        RECT  0.000 195.170 65.000 200.640 ;
        RECT  0.000 201.660 65.000 221.520 ;
        RECT  0.000 222.720 65.000 246.820 ;
        LAYER M2 ;
        RECT  0.000 186.470 65.000 195.650 ;
        LAYER M3 ;
        RECT  64.200 192.330 65.000 200.640 ;
        RECT  0.000 201.660 65.000 221.520 ;
        RECT  0.000 222.720 65.000 246.820 ;
        RECT  0.000 192.330 0.800 200.640 ;
        END
    END VDDO
    PIN VSSO
        DIRECTION INOUT ;
        USE ground ;
        PORT
        LAYER TOP_M ;
        RECT  0.000 92.060 65.000 123.250 ;
        RECT  0.000 155.410 65.000 162.610 ;
        LAYER M2 ;
        RECT  0.000 147.040 65.000 154.520 ;
        LAYER M3 ;
        RECT  0.000 92.060 65.000 123.250 ;
        RECT  64.200 149.940 65.000 162.610 ;
        RECT  0.000 149.940 0.800 162.610 ;
        END
    END VSSO
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        PORT
        LAYER TOP_M ;
        RECT  0.000 123.850 65.000 154.560 ;
        LAYER M2 ;
        RECT  0.000 136.310 65.000 146.340 ;
        LAYER M3 ;
        RECT  64.200 130.690 65.000 148.880 ;
        RECT  0.000 130.690 0.800 148.880 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        PORT
        LAYER TOP_M ;
        RECT  0.000 163.500 65.000 194.560 ;
        LAYER M2 ;
        RECT  0.000 172.080 65.000 183.060 ;
        LAYER M3 ;
        RECT  64.200 163.510 65.000 190.890 ;
        RECT  0.000 163.510 0.800 190.890 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.000 0.000 63.000 250.000 ;
        RECT  0.000 88.990 65.000 130.360 ;
        RECT  0.000 136.510 65.000 157.550 ;
        RECT  0.315 158.150 64.700 158.460 ;
        RECT  0.300 158.930 64.700 159.230 ;
        RECT  0.300 159.530 64.700 159.830 ;
        RECT  0.300 160.130 64.700 160.430 ;
        RECT  0.300 160.730 64.700 161.030 ;
        RECT  0.300 161.330 64.700 161.630 ;
        RECT  0.300 161.910 64.700 162.190 ;
        RECT  0.300 162.490 64.700 162.770 ;
        RECT  0.300 163.070 64.700 163.350 ;
        RECT  0.300 163.650 64.700 163.950 ;
        RECT  0.300 164.250 64.700 164.550 ;
        RECT  0.300 164.850 64.700 165.150 ;
        RECT  0.300 165.450 64.700 165.750 ;
        RECT  0.300 166.050 64.700 166.350 ;
        RECT  0.300 166.650 64.700 166.960 ;
        RECT  0.300 167.260 64.700 167.560 ;
        RECT  0.300 167.860 64.700 168.160 ;
        RECT  0.000 169.150 65.000 197.240 ;
        RECT  0.600 0.600 64.400 250.000 ;
        RECT  0.000 198.470 65.000 250.000 ;
        LAYER M2 ;
        RECT  1.840 196.420 2.120 249.400 ;
        RECT  63.180 196.430 63.670 249.400 ;
        RECT  0.600 196.440 64.400 245.485 ;
        RECT  27.660 196.440 64.400 248.790 ;
        RECT  0.600 196.440 24.080 249.400 ;
        RECT  27.660 196.440 28.080 249.400 ;
        RECT  30.390 196.440 64.400 249.400 ;
        RECT  0.600 183.850 64.400 185.680 ;
        RECT  32.400 155.220 32.720 171.290 ;
        RECT  46.115 155.130 48.355 171.290 ;
        RECT  49.295 155.300 49.605 171.290 ;
        RECT  0.600 155.310 64.400 171.290 ;
        RECT  6.160 155.310 6.440 171.380 ;
        RECT  45.210 155.310 45.490 171.480 ;
        RECT  50.025 155.310 51.995 171.480 ;
        RECT  2.000 0.000 63.000 60.210 ;
        RECT  0.600 0.600 64.400 60.210 ;
        RECT  0.600 0.600 1.210 135.520 ;
        RECT  0.600 91.020 64.400 135.520 ;
        RECT  4.080 91.020 60.940 135.690 ;
        RECT  62.580 91.020 62.995 135.710 ;
        LAYER M3 ;
        RECT  0.600 247.660 24.350 248.740 ;
        RECT  0.600 247.660 24.030 249.400 ;
        RECT  27.390 247.660 64.400 248.740 ;
        RECT  27.710 247.660 28.030 249.400 ;
        RECT  30.440 247.660 64.400 249.400 ;
        RECT  0.600 124.090 64.400 129.850 ;
        RECT  1.640 124.090 63.600 135.790 ;
        RECT  1.810 124.090 2.830 154.520 ;
        RECT  4.040 123.970 60.900 171.560 ;
        RECT  1.640 155.040 63.600 171.560 ;
        RECT  1.640 183.580 63.600 185.950 ;
        RECT  5.490 124.090 63.600 200.820 ;
        RECT  1.640 196.170 63.600 200.820 ;
        RECT  56.930 123.970 57.210 201.060 ;
        RECT  0.600 0.600 64.400 60.480 ;
        RECT  2.000 0.000 63.000 88.700 ;
        RECT  0.600 0.600 1.480 91.220 ;
        RECT  0.600 90.750 64.400 91.220 ;
        LAYER TOP_M ;
        RECT  0.600 247.690 64.400 248.850 ;
        RECT  0.600 247.690 24.140 249.400 ;
        RECT  27.600 247.690 28.140 249.400 ;
        RECT  30.330 247.690 64.400 249.400 ;
        RECT  2.000 0.000 63.000 91.190 ;
        RECT  0.600 0.600 64.400 91.190 ;
    END
END pc3d21d

MACRO pc3d21
    CLASS PAD ;
    FOREIGN pc3d21 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 65.000 BY 250.000 ;
    SYMMETRY X Y R90 ;
    SITE IOSite_c ;
    PIN PAD
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 55.440  LAYER TOP_M  ;
        ANTENNAPARTIALMETALSIDEAREA 287.938  LAYER M3  ;
        ANTENNAPARTIALMETALSIDEAREA 480.740  LAYER M2  ;
        ANTENNADIFFAREA 2657.280  LAYER TOP_M  ;
        ANTENNADIFFAREA 2657.280  LAYER M3  ;
        ANTENNADIFFAREA 1209.600  LAYER M2  ;
        ANTENNAPARTIALCUTAREA 255.798  LAYER V2  ;
        ANTENNAPARTIALCUTAREA 632.318  LAYER TOP_V  ;
        ANTENNAPARTIALCUTAREA 349.898  LAYER V3  ;
        PORT
        LAYER M2 ;
        RECT  2.000 61.000 63.000 90.230 ;
        RECT  24.870 246.275 26.870 250.000 ;
        LAYER M3 ;
        RECT  24.870 249.580 26.870 250.000 ;
        END
    END PAD
    PIN CIN
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 67.374  LAYER M1  ;
        ANTENNAPARTIALMETALSIDEAREA 188.733  LAYER M2  ;
        ANTENNAPARTIALMETALSIDEAREA 40.715  LAYER M3  ;
        ANTENNADIFFAREA 21.020  LAYER M3  ;
        ANTENNADIFFAREA 21.020  LAYER M2  ;
        ANTENNAPARTIALCUTAREA 0.270  LAYER V2  ;
        ANTENNAPARTIALCUTAREA 0.203  LAYER V3  ;
        PORT
        LAYER M2 ;
        RECT  28.870 249.580 29.600 250.000 ;
        LAYER M3 ;
        RECT  28.870 249.580 29.600 250.000 ;
        END
    END CIN
    PIN VDDO
        DIRECTION INOUT ;
        USE power ;
        PORT
        LAYER TOP_M ;
        RECT  0.000 195.170 65.000 200.640 ;
        RECT  0.000 201.660 65.000 221.520 ;
        RECT  0.000 222.720 65.000 246.820 ;
        LAYER M2 ;
        RECT  0.000 186.470 65.000 195.650 ;
        LAYER M3 ;
        RECT  64.200 192.330 65.000 200.640 ;
        RECT  0.000 201.660 65.000 221.520 ;
        RECT  0.000 222.720 65.000 246.820 ;
        RECT  0.000 192.330 0.800 200.640 ;
        END
    END VDDO
    PIN VSSO
        DIRECTION INOUT ;
        USE ground ;
        PORT
        LAYER TOP_M ;
        RECT  0.000 92.060 65.000 123.250 ;
        RECT  0.000 155.410 65.000 162.610 ;
        LAYER M2 ;
        RECT  0.000 147.040 65.000 154.520 ;
        LAYER M3 ;
        RECT  0.000 92.060 65.000 123.250 ;
        RECT  64.200 149.940 65.000 162.610 ;
        RECT  0.000 149.940 0.800 162.610 ;
        END
    END VSSO
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        PORT
        LAYER TOP_M ;
        RECT  0.000 123.850 65.000 154.560 ;
        LAYER M2 ;
        RECT  0.000 136.310 65.000 146.340 ;
        LAYER M3 ;
        RECT  64.200 130.690 65.000 148.880 ;
        RECT  0.000 130.690 0.800 148.880 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        PORT
        LAYER TOP_M ;
        RECT  0.000 163.500 65.000 194.560 ;
        LAYER M2 ;
        RECT  0.000 172.080 65.000 183.060 ;
        LAYER M3 ;
        RECT  64.200 163.510 65.000 190.890 ;
        RECT  0.000 163.510 0.800 190.890 ;
        END
    END VDD
    OBS
        LAYER M1 ;
        RECT  2.000 0.000 63.000 250.000 ;
        RECT  0.000 88.990 65.000 130.360 ;
        RECT  0.000 136.510 65.000 157.550 ;
        RECT  0.315 158.150 64.700 158.460 ;
        RECT  0.300 158.930 64.700 159.230 ;
        RECT  0.300 159.530 64.700 159.830 ;
        RECT  0.300 160.130 64.700 160.430 ;
        RECT  0.300 160.730 64.700 161.030 ;
        RECT  0.300 161.330 64.700 161.630 ;
        RECT  0.300 161.910 64.700 162.190 ;
        RECT  0.300 162.490 64.700 162.770 ;
        RECT  0.300 163.070 64.700 163.350 ;
        RECT  0.300 163.650 64.700 163.950 ;
        RECT  0.300 164.250 64.700 164.550 ;
        RECT  0.300 164.850 64.700 165.150 ;
        RECT  0.300 165.450 64.700 165.750 ;
        RECT  0.300 166.050 64.700 166.350 ;
        RECT  0.300 166.650 64.700 166.960 ;
        RECT  0.300 167.260 64.700 167.560 ;
        RECT  0.300 167.860 64.700 168.160 ;
        RECT  0.000 169.150 65.000 197.240 ;
        RECT  0.600 0.600 64.400 250.000 ;
        RECT  0.000 198.470 65.000 250.000 ;
        LAYER M2 ;
        RECT  1.840 196.420 2.120 249.400 ;
        RECT  63.180 196.430 63.670 249.400 ;
        RECT  0.600 196.440 64.400 245.485 ;
        RECT  27.660 196.440 64.400 248.790 ;
        RECT  0.600 196.440 24.080 249.400 ;
        RECT  27.660 196.440 28.080 249.400 ;
        RECT  30.390 196.440 64.400 249.400 ;
        RECT  0.600 183.850 64.400 185.680 ;
        RECT  32.400 155.220 32.720 171.290 ;
        RECT  0.600 155.310 64.400 171.290 ;
        RECT  6.160 155.310 6.440 171.380 ;
        RECT  45.210 155.310 45.490 171.480 ;
        RECT  50.025 155.310 51.995 171.480 ;
        RECT  2.000 0.000 63.000 60.210 ;
        RECT  0.600 0.600 64.400 60.210 ;
        RECT  0.600 0.600 1.210 135.520 ;
        RECT  0.600 91.020 64.400 135.520 ;
        RECT  4.080 91.020 60.940 135.690 ;
        RECT  62.580 91.020 62.995 135.710 ;
        LAYER M3 ;
        RECT  0.600 247.660 24.350 248.740 ;
        RECT  0.600 247.660 24.030 249.400 ;
        RECT  27.390 247.660 64.400 248.740 ;
        RECT  27.710 247.660 28.030 249.400 ;
        RECT  30.440 247.660 64.400 249.400 ;
        RECT  0.600 124.090 64.400 129.850 ;
        RECT  1.640 124.090 63.600 135.790 ;
        RECT  1.810 124.090 2.830 154.520 ;
        RECT  4.040 123.970 60.900 171.560 ;
        RECT  1.640 155.040 63.600 171.560 ;
        RECT  1.640 183.580 63.600 185.950 ;
        RECT  5.490 124.090 63.600 200.820 ;
        RECT  1.640 196.170 63.600 200.820 ;
        RECT  56.930 123.970 57.210 201.060 ;
        RECT  0.600 0.600 64.400 60.480 ;
        RECT  2.000 0.000 63.000 88.700 ;
        RECT  0.600 0.600 1.480 91.220 ;
        RECT  0.600 90.750 64.400 91.220 ;
        LAYER TOP_M ;
        RECT  0.600 247.690 64.400 248.850 ;
        RECT  0.600 247.690 24.140 249.400 ;
        RECT  27.600 247.690 28.140 249.400 ;
        RECT  30.330 247.690 64.400 249.400 ;
        RECT  2.000 0.000 63.000 91.190 ;
        RECT  0.600 0.600 64.400 91.190 ;
    END
END pc3d21

MACRO pc3d11u
    CLASS PAD ;
    FOREIGN pc3d11u 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 65.000 BY 250.000 ;
    SYMMETRY X Y R90 ;
    SITE IOSite_c ;
    PIN PAD
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 55.440  LAYER TOP_M  ;
        ANTENNAPARTIALMETALSIDEAREA 287.938  LAYER M3  ;
        ANTENNAPARTIALMETALSIDEAREA 480.740  LAYER M2  ;
        ANTENNADIFFAREA 2657.280  LAYER TOP_M  ;
        ANTENNADIFFAREA 2657.280  LAYER M3  ;
        ANTENNADIFFAREA 1209.600  LAYER M2  ;
        ANTENNAPARTIALCUTAREA 255.798  LAYER V2  ;
        ANTENNAPARTIALCUTAREA 632.318  LAYER TOP_V  ;
        ANTENNAPARTIALCUTAREA 349.898  LAYER V3  ;
        PORT
        LAYER M2 ;
        RECT  2.000 61.000 63.000 90.230 ;
        RECT  24.870 246.275 26.870 250.000 ;
        LAYER M3 ;
        RECT  24.870 249.580 26.870 250.000 ;
        END
    END PAD
    PIN CIN
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 67.374  LAYER M1  ;
        ANTENNAPARTIALMETALSIDEAREA 162.710  LAYER M2  ;
        ANTENNAPARTIALMETALSIDEAREA 40.715  LAYER M3  ;
        ANTENNADIFFAREA 3.720  LAYER M2  ;
        ANTENNADIFFAREA 20.600  LAYER M3  ;
        ANTENNAPARTIALCUTAREA 0.203  LAYER V2  ;
        ANTENNAPARTIALCUTAREA 0.203  LAYER V3  ;
        PORT
        LAYER M2 ;
        RECT  28.870 249.580 29.600 250.000 ;
        LAYER M3 ;
        RECT  28.870 249.580 29.600 250.000 ;
        END
    END CIN
    PIN VDDO
        DIRECTION INOUT ;
        USE power ;
        PORT
        LAYER M2 ;
        RECT  0.000 186.470 65.000 195.650 ;
        LAYER M3 ;
        RECT  64.200 192.330 65.000 200.640 ;
        RECT  0.000 201.660 65.000 221.520 ;
        RECT  0.000 222.720 65.000 246.820 ;
        RECT  0.000 192.330 0.800 200.640 ;
        LAYER TOP_M ;
        RECT  0.000 195.170 65.000 200.640 ;
        RECT  0.000 201.660 65.000 221.520 ;
        RECT  0.000 222.720 65.000 246.820 ;
        END
    END VDDO
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        PORT
        LAYER M2 ;
        RECT  0.000 172.080 65.000 183.060 ;
        LAYER M3 ;
        RECT  64.200 163.510 65.000 190.890 ;
        RECT  0.000 163.510 0.800 190.890 ;
        LAYER TOP_M ;
        RECT  0.000 163.500 65.000 194.560 ;
        END
    END VDD
    PIN VSSO
        DIRECTION INOUT ;
        USE ground ;
        PORT
        LAYER M2 ;
        RECT  0.000 147.040 65.000 154.520 ;
        LAYER M3 ;
        RECT  0.000 92.060 65.000 123.250 ;
        RECT  64.200 149.940 65.000 162.610 ;
        RECT  0.000 149.940 0.800 162.610 ;
        LAYER TOP_M ;
        RECT  0.000 92.060 65.000 123.250 ;
        RECT  0.000 155.410 65.000 162.610 ;
        END
    END VSSO
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        PORT
        LAYER M2 ;
        RECT  0.000 136.310 65.000 146.340 ;
        LAYER M3 ;
        RECT  64.200 130.690 65.000 148.880 ;
        RECT  0.000 130.690 0.800 148.880 ;
        LAYER TOP_M ;
        RECT  0.000 123.850 65.000 154.560 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  2.000 0.000 63.000 250.000 ;
        RECT  0.000 88.990 65.000 130.360 ;
        RECT  0.000 136.510 65.000 157.550 ;
        RECT  0.315 158.150 64.700 158.460 ;
        RECT  0.300 158.930 64.700 159.230 ;
        RECT  0.300 159.530 64.700 159.830 ;
        RECT  0.300 160.130 64.700 160.430 ;
        RECT  0.300 160.730 64.700 161.030 ;
        RECT  0.300 161.330 64.700 161.630 ;
        RECT  0.300 161.910 64.700 162.190 ;
        RECT  0.300 162.490 64.700 162.770 ;
        RECT  0.300 163.070 64.700 163.350 ;
        RECT  0.300 163.650 64.700 163.950 ;
        RECT  0.300 164.250 64.700 164.550 ;
        RECT  0.300 164.850 64.700 165.150 ;
        RECT  0.300 165.450 64.700 165.750 ;
        RECT  0.300 166.050 64.700 166.350 ;
        RECT  0.300 166.650 64.700 166.960 ;
        RECT  0.300 167.260 64.700 167.560 ;
        RECT  0.300 167.860 64.700 168.160 ;
        RECT  0.000 169.150 65.000 197.240 ;
        RECT  0.600 0.600 64.400 250.000 ;
        RECT  0.000 198.470 65.000 250.000 ;
        LAYER M2 ;
        RECT  1.840 196.420 2.120 249.400 ;
        RECT  63.180 196.430 63.670 249.400 ;
        RECT  0.600 196.440 64.400 245.485 ;
        RECT  27.660 196.440 64.400 248.790 ;
        RECT  0.600 196.440 24.080 249.400 ;
        RECT  27.660 196.440 28.080 249.400 ;
        RECT  30.390 196.440 64.400 249.400 ;
        RECT  19.440 183.720 30.190 185.680 ;
        RECT  31.430 183.720 52.700 185.680 ;
        RECT  0.600 183.850 64.400 185.680 ;
        RECT  46.260 183.720 51.390 185.710 ;
        RECT  32.450 155.150 32.770 171.290 ;
        RECT  0.600 155.310 64.400 171.290 ;
        RECT  24.770 155.310 25.270 171.375 ;
        RECT  6.160 155.310 6.440 171.380 ;
        RECT  2.000 0.000 63.000 60.210 ;
        RECT  0.600 0.600 64.400 60.210 ;
        RECT  0.600 0.600 1.210 135.520 ;
        RECT  0.600 91.020 64.400 135.520 ;
        RECT  4.080 91.020 60.940 135.690 ;
        RECT  62.580 91.020 62.995 135.710 ;
        LAYER M3 ;
        RECT  0.600 247.660 24.350 248.740 ;
        RECT  0.600 247.660 24.030 249.400 ;
        RECT  27.390 247.660 64.400 248.740 ;
        RECT  27.710 247.660 28.030 249.400 ;
        RECT  30.440 247.660 64.400 249.400 ;
        RECT  0.600 124.090 64.400 129.850 ;
        RECT  1.640 124.090 63.600 135.790 ;
        RECT  1.810 124.090 2.830 154.520 ;
        RECT  4.040 123.970 60.900 171.560 ;
        RECT  1.640 155.040 63.600 171.560 ;
        RECT  1.640 183.580 63.600 185.950 ;
        RECT  5.490 124.090 63.600 200.820 ;
        RECT  1.640 196.170 63.600 200.820 ;
        RECT  56.930 123.970 57.210 201.060 ;
        RECT  0.600 0.600 64.400 60.480 ;
        RECT  2.000 0.000 63.000 88.700 ;
        RECT  0.600 0.600 1.480 91.220 ;
        RECT  0.600 90.750 64.400 91.220 ;
        LAYER TOP_M ;
        RECT  0.600 247.690 64.400 248.850 ;
        RECT  0.600 247.690 24.140 249.400 ;
        RECT  27.600 247.690 28.140 249.400 ;
        RECT  30.330 247.690 64.400 249.400 ;
        RECT  2.000 0.000 63.000 91.190 ;
        RECT  0.600 0.600 64.400 91.190 ;
    END
END pc3d11u

MACRO pc3d11d
    CLASS PAD ;
    FOREIGN pc3d11d 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 65.000 BY 250.000 ;
    SYMMETRY X Y R90 ;
    SITE IOSite_c ;
    PIN PAD
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 55.440  LAYER TOP_M  ;
        ANTENNAPARTIALMETALSIDEAREA 287.938  LAYER M3  ;
        ANTENNAPARTIALMETALSIDEAREA 480.740  LAYER M2  ;
        ANTENNADIFFAREA 2657.280  LAYER TOP_M  ;
        ANTENNADIFFAREA 2657.280  LAYER M3  ;
        ANTENNADIFFAREA 1209.600  LAYER M2  ;
        ANTENNAPARTIALCUTAREA 255.798  LAYER V2  ;
        ANTENNAPARTIALCUTAREA 632.318  LAYER TOP_V  ;
        ANTENNAPARTIALCUTAREA 349.898  LAYER V3  ;
        PORT
        LAYER M2 ;
        RECT  2.000 61.000 63.000 90.230 ;
        RECT  24.870 246.275 26.870 250.000 ;
        LAYER M3 ;
        RECT  24.870 249.580 26.870 250.000 ;
        END
    END PAD
    PIN CIN
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 67.374  LAYER M1  ;
        ANTENNAPARTIALMETALSIDEAREA 162.710  LAYER M2  ;
        ANTENNAPARTIALMETALSIDEAREA 40.715  LAYER M3  ;
        ANTENNADIFFAREA 3.720  LAYER M2  ;
        ANTENNADIFFAREA 20.600  LAYER M3  ;
        ANTENNAPARTIALCUTAREA 0.203  LAYER V2  ;
        ANTENNAPARTIALCUTAREA 0.203  LAYER V3  ;
        PORT
        LAYER M2 ;
        RECT  28.870 249.580 29.600 250.000 ;
        LAYER M3 ;
        RECT  28.870 249.580 29.600 250.000 ;
        END
    END CIN
    PIN VDDO
        DIRECTION INOUT ;
        USE power ;
        PORT
        LAYER M2 ;
        RECT  0.000 186.470 65.000 195.650 ;
        LAYER M3 ;
        RECT  64.200 192.330 65.000 200.640 ;
        RECT  0.000 201.660 65.000 221.520 ;
        RECT  0.000 222.720 65.000 246.820 ;
        RECT  0.000 192.330 0.800 200.640 ;
        LAYER TOP_M ;
        RECT  0.000 195.170 65.000 200.640 ;
        RECT  0.000 201.660 65.000 221.520 ;
        RECT  0.000 222.720 65.000 246.820 ;
        END
    END VDDO
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        PORT
        LAYER M2 ;
        RECT  0.000 172.080 65.000 183.060 ;
        LAYER M3 ;
        RECT  64.200 163.510 65.000 190.890 ;
        RECT  0.000 163.510 0.800 190.890 ;
        LAYER TOP_M ;
        RECT  0.000 163.500 65.000 194.560 ;
        END
    END VDD
    PIN VSSO
        DIRECTION INOUT ;
        USE ground ;
        PORT
        LAYER M2 ;
        RECT  0.000 147.040 65.000 154.520 ;
        LAYER M3 ;
        RECT  0.000 92.060 65.000 123.250 ;
        RECT  64.200 149.940 65.000 162.610 ;
        RECT  0.000 149.940 0.800 162.610 ;
        LAYER TOP_M ;
        RECT  0.000 92.060 65.000 123.250 ;
        RECT  0.000 155.410 65.000 162.610 ;
        END
    END VSSO
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        PORT
        LAYER M2 ;
        RECT  0.000 136.310 65.000 146.340 ;
        LAYER M3 ;
        RECT  64.200 130.690 65.000 148.880 ;
        RECT  0.000 130.690 0.800 148.880 ;
        LAYER TOP_M ;
        RECT  0.000 123.850 65.000 154.560 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  2.000 0.000 63.000 250.000 ;
        RECT  0.000 88.990 65.000 130.360 ;
        RECT  0.000 136.510 65.000 157.550 ;
        RECT  0.315 158.150 64.700 158.460 ;
        RECT  0.300 158.930 64.700 159.230 ;
        RECT  0.300 159.530 64.700 159.830 ;
        RECT  0.300 160.130 64.700 160.430 ;
        RECT  0.300 160.730 64.700 161.030 ;
        RECT  0.300 161.330 64.700 161.630 ;
        RECT  0.300 161.910 64.700 162.190 ;
        RECT  0.300 162.490 64.700 162.770 ;
        RECT  0.300 163.070 64.700 163.350 ;
        RECT  0.300 163.650 64.700 163.950 ;
        RECT  0.300 164.250 64.700 164.550 ;
        RECT  0.300 164.850 64.700 165.150 ;
        RECT  0.300 165.450 64.700 165.750 ;
        RECT  0.300 166.050 64.700 166.350 ;
        RECT  0.300 166.650 64.700 166.960 ;
        RECT  0.300 167.260 64.700 167.560 ;
        RECT  0.300 167.860 64.700 168.160 ;
        RECT  0.000 169.150 65.000 197.240 ;
        RECT  0.600 0.600 64.400 250.000 ;
        RECT  0.000 198.470 65.000 250.000 ;
        LAYER M2 ;
        RECT  1.840 196.420 2.120 249.400 ;
        RECT  63.180 196.430 63.670 249.400 ;
        RECT  0.600 196.440 64.400 245.485 ;
        RECT  27.660 196.440 64.400 248.790 ;
        RECT  0.600 196.440 24.080 249.400 ;
        RECT  27.660 196.440 28.080 249.400 ;
        RECT  30.390 196.440 64.400 249.400 ;
        RECT  19.440 183.720 30.190 185.680 ;
        RECT  31.430 183.720 52.700 185.680 ;
        RECT  0.600 183.850 64.400 185.680 ;
        RECT  46.260 183.720 51.390 185.710 ;
        RECT  32.450 155.150 32.770 171.290 ;
        RECT  53.030 155.130 55.270 171.290 ;
        RECT  56.210 155.300 56.520 171.290 ;
        RECT  0.600 155.310 64.400 171.290 ;
        RECT  6.160 155.310 6.440 171.380 ;
        RECT  2.000 0.000 63.000 60.210 ;
        RECT  0.600 0.600 64.400 60.210 ;
        RECT  0.600 0.600 1.210 135.520 ;
        RECT  0.600 91.020 64.400 135.520 ;
        RECT  4.080 91.020 60.940 135.690 ;
        RECT  62.580 91.020 62.995 135.710 ;
        LAYER M3 ;
        RECT  0.600 247.660 24.350 248.740 ;
        RECT  0.600 247.660 24.030 249.400 ;
        RECT  27.390 247.660 64.400 248.740 ;
        RECT  27.710 247.660 28.030 249.400 ;
        RECT  30.440 247.660 64.400 249.400 ;
        RECT  0.600 124.090 64.400 129.850 ;
        RECT  1.640 124.090 63.600 135.790 ;
        RECT  1.810 124.090 2.830 154.520 ;
        RECT  4.040 123.970 60.900 171.560 ;
        RECT  1.640 155.040 63.600 171.560 ;
        RECT  1.640 183.580 63.600 185.950 ;
        RECT  5.490 124.090 63.600 200.820 ;
        RECT  1.640 196.170 63.600 200.820 ;
        RECT  56.930 123.970 57.210 201.060 ;
        RECT  0.600 0.600 64.400 60.480 ;
        RECT  2.000 0.000 63.000 88.700 ;
        RECT  0.600 0.600 1.480 91.220 ;
        RECT  0.600 90.750 64.400 91.220 ;
        LAYER TOP_M ;
        RECT  0.600 247.690 64.400 248.850 ;
        RECT  0.600 247.690 24.140 249.400 ;
        RECT  27.600 247.690 28.140 249.400 ;
        RECT  30.330 247.690 64.400 249.400 ;
        RECT  2.000 0.000 63.000 91.190 ;
        RECT  0.600 0.600 64.400 91.190 ;
    END
END pc3d11d

MACRO pc3d11
    CLASS PAD ;
    FOREIGN pc3d11 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 65.000 BY 250.000 ;
    SYMMETRY X Y R90 ;
    SITE IOSite_c ;
    PIN PAD
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 55.440  LAYER TOP_M  ;
        ANTENNAPARTIALMETALSIDEAREA 287.938  LAYER M3  ;
        ANTENNAPARTIALMETALSIDEAREA 480.740  LAYER M2  ;
        ANTENNADIFFAREA 2657.280  LAYER TOP_M  ;
        ANTENNADIFFAREA 2657.280  LAYER M3  ;
        ANTENNADIFFAREA 1209.600  LAYER M2  ;
        ANTENNAPARTIALCUTAREA 255.798  LAYER V2  ;
        ANTENNAPARTIALCUTAREA 632.318  LAYER TOP_V  ;
        ANTENNAPARTIALCUTAREA 349.898  LAYER V3  ;
        PORT
        LAYER M2 ;
        RECT  2.000 61.000 63.000 90.230 ;
        RECT  24.870 246.275 26.870 250.000 ;
        LAYER M3 ;
        RECT  24.870 249.580 26.870 250.000 ;
        END
    END PAD
    PIN CIN
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 67.374  LAYER M1  ;
        ANTENNAPARTIALMETALSIDEAREA 162.710  LAYER M2  ;
        ANTENNAPARTIALMETALSIDEAREA 40.715  LAYER M3  ;
        ANTENNADIFFAREA 3.720  LAYER M2  ;
        ANTENNADIFFAREA 20.600  LAYER M3  ;
        ANTENNAPARTIALCUTAREA 0.203  LAYER V2  ;
        ANTENNAPARTIALCUTAREA 0.203  LAYER V3  ;
        PORT
        LAYER M2 ;
        RECT  28.870 249.580 29.600 250.000 ;
        LAYER M3 ;
        RECT  28.870 249.580 29.600 250.000 ;
        END
    END CIN
    PIN VDDO
        DIRECTION INOUT ;
        USE power ;
        PORT
        LAYER M2 ;
        RECT  0.000 186.470 65.000 195.650 ;
        LAYER M3 ;
        RECT  64.200 192.330 65.000 200.640 ;
        RECT  0.000 201.660 65.000 221.520 ;
        RECT  0.000 222.720 65.000 246.820 ;
        RECT  0.000 192.330 0.800 200.640 ;
        LAYER TOP_M ;
        RECT  0.000 195.170 65.000 200.640 ;
        RECT  0.000 201.660 65.000 221.520 ;
        RECT  0.000 222.720 65.000 246.820 ;
        END
    END VDDO
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        PORT
        LAYER M2 ;
        RECT  0.000 172.080 65.000 183.060 ;
        LAYER M3 ;
        RECT  64.200 163.510 65.000 190.890 ;
        RECT  0.000 163.510 0.800 190.890 ;
        LAYER TOP_M ;
        RECT  0.000 163.500 65.000 194.560 ;
        END
    END VDD
    PIN VSSO
        DIRECTION INOUT ;
        USE ground ;
        PORT
        LAYER M2 ;
        RECT  0.000 147.040 65.000 154.520 ;
        LAYER M3 ;
        RECT  0.000 92.060 65.000 123.250 ;
        RECT  64.200 149.940 65.000 162.610 ;
        RECT  0.000 149.940 0.800 162.610 ;
        LAYER TOP_M ;
        RECT  0.000 92.060 65.000 123.250 ;
        RECT  0.000 155.410 65.000 162.610 ;
        END
    END VSSO
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        PORT
        LAYER M2 ;
        RECT  0.000 136.310 65.000 146.340 ;
        LAYER M3 ;
        RECT  64.200 130.690 65.000 148.880 ;
        RECT  0.000 130.690 0.800 148.880 ;
        LAYER TOP_M ;
        RECT  0.000 123.850 65.000 154.560 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  2.000 0.000 63.000 250.000 ;
        RECT  0.000 88.990 65.000 130.360 ;
        RECT  0.000 136.510 65.000 157.550 ;
        RECT  0.315 158.150 64.700 158.460 ;
        RECT  0.300 158.930 64.700 159.230 ;
        RECT  0.300 159.530 64.700 159.830 ;
        RECT  0.300 160.130 64.700 160.430 ;
        RECT  0.300 160.730 64.700 161.030 ;
        RECT  0.300 161.330 64.700 161.630 ;
        RECT  0.300 161.910 64.700 162.190 ;
        RECT  0.300 162.490 64.700 162.770 ;
        RECT  0.300 163.070 64.700 163.350 ;
        RECT  0.300 163.650 64.700 163.950 ;
        RECT  0.300 164.250 64.700 164.550 ;
        RECT  0.300 164.850 64.700 165.150 ;
        RECT  0.300 165.450 64.700 165.750 ;
        RECT  0.300 166.050 64.700 166.350 ;
        RECT  0.300 166.650 64.700 166.960 ;
        RECT  0.300 167.260 64.700 167.560 ;
        RECT  0.300 167.860 64.700 168.160 ;
        RECT  0.000 169.150 65.000 197.240 ;
        RECT  0.600 0.600 64.400 250.000 ;
        RECT  0.000 198.470 65.000 250.000 ;
        LAYER M2 ;
        RECT  1.840 196.420 2.120 249.400 ;
        RECT  63.180 196.430 63.670 249.400 ;
        RECT  0.600 196.440 64.400 245.485 ;
        RECT  27.660 196.440 64.400 248.790 ;
        RECT  0.600 196.440 24.080 249.400 ;
        RECT  27.660 196.440 28.080 249.400 ;
        RECT  30.390 196.440 64.400 249.400 ;
        RECT  19.440 183.720 30.190 185.680 ;
        RECT  31.430 183.720 52.700 185.680 ;
        RECT  0.600 183.850 64.400 185.680 ;
        RECT  46.260 183.720 51.390 185.710 ;
        RECT  32.450 155.150 32.770 171.290 ;
        RECT  0.600 155.310 64.400 171.290 ;
        RECT  6.160 155.310 6.440 171.380 ;
        RECT  2.000 0.000 63.000 60.210 ;
        RECT  0.600 0.600 64.400 60.210 ;
        RECT  0.600 0.600 1.210 135.520 ;
        RECT  0.600 91.020 64.400 135.520 ;
        RECT  4.080 91.020 60.940 135.690 ;
        RECT  62.580 91.020 62.995 135.710 ;
        LAYER M3 ;
        RECT  0.600 247.660 24.350 248.740 ;
        RECT  0.600 247.660 24.030 249.400 ;
        RECT  27.390 247.660 64.400 248.740 ;
        RECT  27.710 247.660 28.030 249.400 ;
        RECT  30.440 247.660 64.400 249.400 ;
        RECT  0.600 124.090 64.400 129.850 ;
        RECT  1.640 124.090 63.600 135.790 ;
        RECT  1.810 124.090 2.830 154.520 ;
        RECT  4.040 123.970 60.900 171.560 ;
        RECT  1.640 155.040 63.600 171.560 ;
        RECT  1.640 183.580 63.600 185.950 ;
        RECT  5.490 124.090 63.600 200.820 ;
        RECT  1.640 196.170 63.600 200.820 ;
        RECT  56.930 123.970 57.210 201.060 ;
        RECT  0.600 0.600 64.400 60.480 ;
        RECT  2.000 0.000 63.000 88.700 ;
        RECT  0.600 0.600 1.480 91.220 ;
        RECT  0.600 90.750 64.400 91.220 ;
        LAYER TOP_M ;
        RECT  0.600 247.690 64.400 248.850 ;
        RECT  0.600 247.690 24.140 249.400 ;
        RECT  27.600 247.690 28.140 249.400 ;
        RECT  30.330 247.690 64.400 249.400 ;
        RECT  2.000 0.000 63.000 91.190 ;
        RECT  0.600 0.600 64.400 91.190 ;
    END
END pc3d11

MACRO pc3d01u
    CLASS PAD ;
    FOREIGN pc3d01u 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 65.000 BY 250.000 ;
    SYMMETRY X Y R90 ;
    SITE IOSite_c ;
    PIN PAD
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 55.440  LAYER TOP_M  ;
        ANTENNAPARTIALMETALSIDEAREA 287.938  LAYER M3  ;
        ANTENNAPARTIALMETALSIDEAREA 480.740  LAYER M2  ;
        ANTENNADIFFAREA 2657.280  LAYER TOP_M  ;
        ANTENNADIFFAREA 2657.280  LAYER M3  ;
        ANTENNADIFFAREA 1209.600  LAYER M2  ;
        ANTENNAPARTIALCUTAREA 632.318  LAYER TOP_V  ;
        ANTENNAPARTIALCUTAREA 349.898  LAYER V3  ;
        ANTENNAPARTIALCUTAREA 255.798  LAYER V2  ;
        PORT
        LAYER M2 ;
        RECT  2.000 61.000 63.000 90.230 ;
        RECT  24.870 246.275 26.870 250.000 ;
        LAYER M3 ;
        RECT  24.870 249.580 26.870 250.000 ;
        END
    END PAD
    PIN CIN
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 67.374  LAYER M1  ;
        ANTENNAPARTIALMETALSIDEAREA 162.668  LAYER M2  ;
        ANTENNAPARTIALMETALSIDEAREA 40.715  LAYER M3  ;
        ANTENNADIFFAREA 3.720  LAYER M2  ;
        ANTENNADIFFAREA 20.600  LAYER M3  ;
        ANTENNAPARTIALCUTAREA 0.203  LAYER V2  ;
        ANTENNAPARTIALCUTAREA 0.203  LAYER V3  ;
        PORT
        LAYER M2 ;
        RECT  28.870 249.580 29.600 250.000 ;
        LAYER M3 ;
        RECT  28.870 249.580 29.600 250.000 ;
        END
    END CIN
    PIN VDDO
        DIRECTION INOUT ;
        USE power ;
        PORT
        LAYER M2 ;
        RECT  0.000 186.470 65.000 195.650 ;
        LAYER M3 ;
        RECT  64.200 192.330 65.000 200.640 ;
        RECT  0.000 201.660 65.000 221.520 ;
        RECT  0.000 222.720 65.000 246.820 ;
        RECT  0.000 192.330 0.800 200.640 ;
        LAYER TOP_M ;
        RECT  0.000 195.170 65.000 200.640 ;
        RECT  0.000 201.660 65.000 221.520 ;
        RECT  0.000 222.720 65.000 246.820 ;
        END
    END VDDO
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        PORT
        LAYER M2 ;
        RECT  0.000 172.080 65.000 183.060 ;
        LAYER M3 ;
        RECT  64.200 163.510 65.000 190.890 ;
        RECT  0.000 163.510 0.800 190.890 ;
        LAYER TOP_M ;
        RECT  0.000 163.500 65.000 194.560 ;
        END
    END VDD
    PIN VSSO
        DIRECTION INOUT ;
        USE ground ;
        PORT
        LAYER M2 ;
        RECT  0.000 147.040 65.000 154.520 ;
        LAYER M3 ;
        RECT  0.000 92.060 65.000 123.250 ;
        RECT  64.200 149.940 65.000 162.610 ;
        RECT  0.000 149.940 0.800 162.610 ;
        LAYER TOP_M ;
        RECT  0.000 92.060 65.000 123.250 ;
        RECT  0.000 155.410 65.000 162.610 ;
        END
    END VSSO
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        PORT
        LAYER M2 ;
        RECT  0.000 136.310 65.000 146.340 ;
        LAYER M3 ;
        RECT  64.200 130.690 65.000 148.880 ;
        RECT  0.000 130.690 0.800 148.880 ;
        LAYER TOP_M ;
        RECT  0.000 123.850 65.000 154.560 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  2.000 0.000 63.000 250.000 ;
        RECT  0.000 88.990 65.000 130.360 ;
        RECT  0.000 136.510 65.000 157.550 ;
        RECT  0.315 158.150 64.700 158.460 ;
        RECT  0.300 158.930 64.700 159.230 ;
        RECT  0.300 159.530 64.700 159.830 ;
        RECT  0.300 160.130 64.700 160.430 ;
        RECT  0.300 160.730 64.700 161.030 ;
        RECT  0.300 161.330 64.700 161.630 ;
        RECT  0.300 161.910 64.700 162.190 ;
        RECT  0.300 162.490 64.700 162.770 ;
        RECT  0.300 163.070 64.700 163.350 ;
        RECT  0.300 163.650 64.700 163.950 ;
        RECT  0.300 164.250 64.700 164.550 ;
        RECT  0.300 164.850 64.700 165.150 ;
        RECT  0.300 165.450 64.700 165.750 ;
        RECT  0.300 166.050 64.700 166.350 ;
        RECT  0.300 166.650 64.700 166.960 ;
        RECT  0.300 167.260 64.700 167.560 ;
        RECT  0.300 167.860 64.700 168.160 ;
        RECT  0.000 169.150 65.000 197.240 ;
        RECT  0.600 0.600 64.400 250.000 ;
        RECT  0.000 198.470 65.000 250.000 ;
        LAYER M2 ;
        RECT  1.840 196.420 2.120 249.400 ;
        RECT  63.180 196.430 63.670 249.400 ;
        RECT  0.600 196.440 64.400 245.485 ;
        RECT  27.660 196.440 64.400 248.790 ;
        RECT  0.600 196.440 24.080 249.400 ;
        RECT  27.660 196.440 28.080 249.400 ;
        RECT  30.390 196.440 64.400 249.400 ;
        RECT  19.440 183.720 52.270 185.680 ;
        RECT  0.600 183.850 64.400 185.680 ;
        RECT  46.260 183.720 51.390 185.710 ;
        RECT  0.600 155.310 64.400 171.290 ;
        RECT  24.710 155.310 25.210 171.375 ;
        RECT  6.160 155.310 6.440 171.380 ;
        RECT  2.000 0.000 63.000 60.210 ;
        RECT  0.600 0.600 64.400 60.210 ;
        RECT  0.600 0.600 1.210 135.520 ;
        RECT  0.600 91.020 64.400 135.520 ;
        RECT  4.080 91.020 60.940 135.690 ;
        RECT  62.580 91.020 62.995 135.710 ;
        LAYER M3 ;
        RECT  0.600 247.660 24.350 248.740 ;
        RECT  0.600 247.660 24.030 249.400 ;
        RECT  27.390 247.660 64.400 248.740 ;
        RECT  27.710 247.660 28.030 249.400 ;
        RECT  30.440 247.660 64.400 249.400 ;
        RECT  0.600 124.090 64.400 129.850 ;
        RECT  1.640 124.090 63.600 135.790 ;
        RECT  1.810 124.090 2.830 154.520 ;
        RECT  4.040 123.970 60.900 171.560 ;
        RECT  1.640 155.040 63.600 171.560 ;
        RECT  1.640 183.580 63.600 185.950 ;
        RECT  5.490 124.090 63.600 200.820 ;
        RECT  1.640 196.170 63.600 200.820 ;
        RECT  56.930 123.970 57.210 201.060 ;
        RECT  0.600 0.600 64.400 60.480 ;
        RECT  2.000 0.000 63.000 88.700 ;
        RECT  0.600 0.600 1.480 91.220 ;
        RECT  0.600 90.750 64.400 91.220 ;
        LAYER TOP_M ;
        RECT  0.600 247.690 64.400 248.850 ;
        RECT  0.600 247.690 24.140 249.400 ;
        RECT  27.600 247.690 28.140 249.400 ;
        RECT  30.330 247.690 64.400 249.400 ;
        RECT  2.000 0.000 63.000 91.190 ;
        RECT  0.600 0.600 64.400 91.190 ;
    END
END pc3d01u

MACRO pc3d01d
    CLASS PAD ;
    FOREIGN pc3d01d 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 65.000 BY 250.000 ;
    SYMMETRY X Y R90 ;
    SITE IOSite_c ;
    PIN PAD
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 55.440  LAYER TOP_M  ;
        ANTENNAPARTIALMETALSIDEAREA 287.938  LAYER M3  ;
        ANTENNAPARTIALMETALSIDEAREA 480.740  LAYER M2  ;
        ANTENNADIFFAREA 2657.280  LAYER TOP_M  ;
        ANTENNADIFFAREA 2657.280  LAYER M3  ;
        ANTENNADIFFAREA 1209.600  LAYER M2  ;
        ANTENNAPARTIALCUTAREA 632.318  LAYER TOP_V  ;
        ANTENNAPARTIALCUTAREA 349.898  LAYER V3  ;
        ANTENNAPARTIALCUTAREA 255.798  LAYER V2  ;
        PORT
        LAYER M2 ;
        RECT  2.000 61.000 63.000 90.230 ;
        RECT  24.870 246.275 26.870 250.000 ;
        LAYER M3 ;
        RECT  24.870 249.580 26.870 250.000 ;
        END
    END PAD
    PIN CIN
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 67.374  LAYER M1  ;
        ANTENNAPARTIALMETALSIDEAREA 162.668  LAYER M2  ;
        ANTENNAPARTIALMETALSIDEAREA 40.715  LAYER M3  ;
        ANTENNADIFFAREA 3.720  LAYER M2  ;
        ANTENNADIFFAREA 20.600  LAYER M3  ;
        ANTENNAPARTIALCUTAREA 0.203  LAYER V2  ;
        ANTENNAPARTIALCUTAREA 0.203  LAYER V3  ;
        PORT
        LAYER M2 ;
        RECT  28.870 249.580 29.600 250.000 ;
        LAYER M3 ;
        RECT  28.870 249.580 29.600 250.000 ;
        END
    END CIN
    PIN VDDO
        DIRECTION INOUT ;
        USE power ;
        PORT
        LAYER M2 ;
        RECT  0.000 186.470 65.000 195.650 ;
        LAYER M3 ;
        RECT  64.200 192.330 65.000 200.640 ;
        RECT  0.000 201.660 65.000 221.520 ;
        RECT  0.000 222.720 65.000 246.820 ;
        RECT  0.000 192.330 0.800 200.640 ;
        LAYER TOP_M ;
        RECT  0.000 195.170 65.000 200.640 ;
        RECT  0.000 201.660 65.000 221.520 ;
        RECT  0.000 222.720 65.000 246.820 ;
        END
    END VDDO
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        PORT
        LAYER M2 ;
        RECT  0.000 172.080 65.000 183.060 ;
        LAYER M3 ;
        RECT  64.200 163.510 65.000 190.890 ;
        RECT  0.000 163.510 0.800 190.890 ;
        LAYER TOP_M ;
        RECT  0.000 163.500 65.000 194.560 ;
        END
    END VDD
    PIN VSSO
        DIRECTION INOUT ;
        USE ground ;
        PORT
        LAYER M2 ;
        RECT  0.000 147.040 65.000 154.520 ;
        LAYER M3 ;
        RECT  0.000 92.060 65.000 123.250 ;
        RECT  64.200 149.940 65.000 162.610 ;
        RECT  0.000 149.940 0.800 162.610 ;
        LAYER TOP_M ;
        RECT  0.000 92.060 65.000 123.250 ;
        RECT  0.000 155.410 65.000 162.610 ;
        END
    END VSSO
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        PORT
        LAYER M2 ;
        RECT  0.000 136.310 65.000 146.340 ;
        LAYER M3 ;
        RECT  64.200 130.690 65.000 148.880 ;
        RECT  0.000 130.690 0.800 148.880 ;
        LAYER TOP_M ;
        RECT  0.000 123.850 65.000 154.560 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  2.000 0.000 63.000 250.000 ;
        RECT  0.000 88.990 65.000 130.360 ;
        RECT  0.000 136.510 65.000 157.550 ;
        RECT  0.315 158.150 64.700 158.460 ;
        RECT  0.300 158.930 64.700 159.230 ;
        RECT  0.300 159.530 64.700 159.830 ;
        RECT  0.300 160.130 64.700 160.430 ;
        RECT  0.300 160.730 64.700 161.030 ;
        RECT  0.300 161.330 64.700 161.630 ;
        RECT  0.300 161.910 64.700 162.190 ;
        RECT  0.300 162.490 64.700 162.770 ;
        RECT  0.300 163.070 64.700 163.350 ;
        RECT  0.300 163.650 64.700 163.950 ;
        RECT  0.300 164.250 64.700 164.550 ;
        RECT  0.300 164.850 64.700 165.150 ;
        RECT  0.300 165.450 64.700 165.750 ;
        RECT  0.300 166.050 64.700 166.350 ;
        RECT  0.300 166.650 64.700 166.960 ;
        RECT  0.300 167.260 64.700 167.560 ;
        RECT  0.300 167.860 64.700 168.160 ;
        RECT  0.000 169.150 65.000 197.240 ;
        RECT  0.600 0.600 64.400 250.000 ;
        RECT  0.000 198.470 65.000 250.000 ;
        LAYER M2 ;
        RECT  1.840 196.420 2.120 249.400 ;
        RECT  63.180 196.430 63.670 249.400 ;
        RECT  0.600 196.440 64.400 245.485 ;
        RECT  27.660 196.440 64.400 248.790 ;
        RECT  0.600 196.440 24.080 249.400 ;
        RECT  27.660 196.440 28.080 249.400 ;
        RECT  30.390 196.440 64.400 249.400 ;
        RECT  19.440 183.720 52.270 185.680 ;
        RECT  0.600 183.850 64.400 185.680 ;
        RECT  46.260 183.720 51.390 185.710 ;
        RECT  44.665 155.130 46.905 171.290 ;
        RECT  47.845 155.300 48.155 171.290 ;
        RECT  0.600 155.310 64.400 171.290 ;
        RECT  6.160 155.310 6.440 171.380 ;
        RECT  2.000 0.000 63.000 60.210 ;
        RECT  0.600 0.600 64.400 60.210 ;
        RECT  0.600 0.600 1.210 135.520 ;
        RECT  0.600 91.020 64.400 135.520 ;
        RECT  4.080 91.020 60.940 135.690 ;
        RECT  62.580 91.020 62.995 135.710 ;
        LAYER M3 ;
        RECT  0.600 247.660 24.350 248.740 ;
        RECT  0.600 247.660 24.030 249.400 ;
        RECT  27.390 247.660 64.400 248.740 ;
        RECT  27.710 247.660 28.030 249.400 ;
        RECT  30.440 247.660 64.400 249.400 ;
        RECT  0.600 124.090 64.400 129.850 ;
        RECT  1.640 124.090 63.600 135.790 ;
        RECT  1.810 124.090 2.830 154.520 ;
        RECT  4.040 123.970 60.900 171.560 ;
        RECT  1.640 155.040 63.600 171.560 ;
        RECT  1.640 183.580 63.600 185.950 ;
        RECT  5.490 124.090 63.600 200.820 ;
        RECT  1.640 196.170 63.600 200.820 ;
        RECT  56.930 123.970 57.210 201.060 ;
        RECT  0.600 0.600 64.400 60.480 ;
        RECT  2.000 0.000 63.000 88.700 ;
        RECT  0.600 0.600 1.480 91.220 ;
        RECT  0.600 90.750 64.400 91.220 ;
        LAYER TOP_M ;
        RECT  0.600 247.690 64.400 248.850 ;
        RECT  0.600 247.690 24.140 249.400 ;
        RECT  27.600 247.690 28.140 249.400 ;
        RECT  30.330 247.690 64.400 249.400 ;
        RECT  2.000 0.000 63.000 91.190 ;
        RECT  0.600 0.600 64.400 91.190 ;
    END
END pc3d01d

MACRO pc3d01
    CLASS PAD ;
    FOREIGN pc3d01 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 65.000 BY 250.000 ;
    SYMMETRY X Y R90 ;
    SITE IOSite_c ;
    PIN PAD
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 55.440  LAYER TOP_M  ;
        ANTENNAPARTIALMETALSIDEAREA 287.938  LAYER M3  ;
        ANTENNAPARTIALMETALSIDEAREA 480.740  LAYER M2  ;
        ANTENNADIFFAREA 2657.280  LAYER TOP_M  ;
        ANTENNADIFFAREA 2657.280  LAYER M3  ;
        ANTENNADIFFAREA 1209.600  LAYER M2  ;
        ANTENNAPARTIALCUTAREA 632.318  LAYER TOP_V  ;
        ANTENNAPARTIALCUTAREA 349.898  LAYER V3  ;
        ANTENNAPARTIALCUTAREA 255.798  LAYER V2  ;
        PORT
        LAYER M2 ;
        RECT  2.000 61.000 63.000 90.230 ;
        RECT  24.870 246.275 26.870 250.000 ;
        LAYER M3 ;
        RECT  24.870 249.580 26.870 250.000 ;
        END
    END PAD
    PIN CIN
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 67.374  LAYER M1  ;
        ANTENNAPARTIALMETALSIDEAREA 162.668  LAYER M2  ;
        ANTENNAPARTIALMETALSIDEAREA 40.715  LAYER M3  ;
        ANTENNADIFFAREA 3.720  LAYER M2  ;
        ANTENNADIFFAREA 20.600  LAYER M3  ;
        ANTENNAPARTIALCUTAREA 0.203  LAYER V2  ;
        ANTENNAPARTIALCUTAREA 0.203  LAYER V3  ;
        PORT
        LAYER M2 ;
        RECT  28.870 249.580 29.600 250.000 ;
        LAYER M3 ;
        RECT  28.870 249.580 29.600 250.000 ;
        END
    END CIN
    PIN VDDO
        DIRECTION INOUT ;
        USE power ;
        PORT
        LAYER M2 ;
        RECT  0.000 186.470 65.000 195.650 ;
        LAYER M3 ;
        RECT  64.200 192.330 65.000 200.640 ;
        RECT  0.000 201.660 65.000 221.520 ;
        RECT  0.000 222.720 65.000 246.820 ;
        RECT  0.000 192.330 0.800 200.640 ;
        LAYER TOP_M ;
        RECT  0.000 195.170 65.000 200.640 ;
        RECT  0.000 201.660 65.000 221.520 ;
        RECT  0.000 222.720 65.000 246.820 ;
        END
    END VDDO
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        PORT
        LAYER M2 ;
        RECT  0.000 172.080 65.000 183.060 ;
        LAYER M3 ;
        RECT  64.200 163.510 65.000 190.890 ;
        RECT  0.000 163.510 0.800 190.890 ;
        LAYER TOP_M ;
        RECT  0.000 163.500 65.000 194.560 ;
        END
    END VDD
    PIN VSSO
        DIRECTION INOUT ;
        USE ground ;
        PORT
        LAYER M2 ;
        RECT  0.000 147.040 65.000 154.520 ;
        LAYER M3 ;
        RECT  0.000 92.060 65.000 123.250 ;
        RECT  64.200 149.940 65.000 162.610 ;
        RECT  0.000 149.940 0.800 162.610 ;
        LAYER TOP_M ;
        RECT  0.000 92.060 65.000 123.250 ;
        RECT  0.000 155.410 65.000 162.610 ;
        END
    END VSSO
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        PORT
        LAYER M2 ;
        RECT  0.000 136.310 65.000 146.340 ;
        LAYER M3 ;
        RECT  64.200 130.690 65.000 148.880 ;
        RECT  0.000 130.690 0.800 148.880 ;
        LAYER TOP_M ;
        RECT  0.000 123.850 65.000 154.560 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  2.000 0.000 63.000 250.000 ;
        RECT  0.000 88.990 65.000 130.360 ;
        RECT  0.000 136.510 65.000 157.550 ;
        RECT  0.315 158.150 64.700 158.460 ;
        RECT  0.300 158.930 64.700 159.230 ;
        RECT  0.300 159.530 64.700 159.830 ;
        RECT  0.300 160.130 64.700 160.430 ;
        RECT  0.300 160.730 64.700 161.030 ;
        RECT  0.300 161.330 64.700 161.630 ;
        RECT  0.300 161.910 64.700 162.190 ;
        RECT  0.300 162.490 64.700 162.770 ;
        RECT  0.300 163.070 64.700 163.350 ;
        RECT  0.300 163.650 64.700 163.950 ;
        RECT  0.300 164.250 64.700 164.550 ;
        RECT  0.300 164.850 64.700 165.150 ;
        RECT  0.300 165.450 64.700 165.750 ;
        RECT  0.300 166.050 64.700 166.350 ;
        RECT  0.300 166.650 64.700 166.960 ;
        RECT  0.300 167.260 64.700 167.560 ;
        RECT  0.300 167.860 64.700 168.160 ;
        RECT  0.000 169.150 65.000 197.240 ;
        RECT  0.600 0.600 64.400 250.000 ;
        RECT  0.000 198.470 65.000 250.000 ;
        LAYER M2 ;
        RECT  1.840 196.420 2.120 249.400 ;
        RECT  63.180 196.430 63.670 249.400 ;
        RECT  0.600 196.440 64.400 245.485 ;
        RECT  27.660 196.440 64.400 248.790 ;
        RECT  0.600 196.440 24.080 249.400 ;
        RECT  27.660 196.440 28.080 249.400 ;
        RECT  30.390 196.440 64.400 249.400 ;
        RECT  19.440 183.720 52.270 185.680 ;
        RECT  0.600 183.850 64.400 185.680 ;
        RECT  46.260 183.720 51.390 185.710 ;
        RECT  0.600 155.310 64.400 171.290 ;
        RECT  6.160 155.310 6.440 171.380 ;
        RECT  2.000 0.000 63.000 60.210 ;
        RECT  0.600 0.600 64.400 60.210 ;
        RECT  0.600 0.600 1.210 135.520 ;
        RECT  0.600 91.020 64.400 135.520 ;
        RECT  4.080 91.020 60.940 135.690 ;
        RECT  62.580 91.020 62.995 135.710 ;
        LAYER M3 ;
        RECT  0.600 247.660 24.350 248.740 ;
        RECT  0.600 247.660 24.030 249.400 ;
        RECT  27.390 247.660 64.400 248.740 ;
        RECT  27.710 247.660 28.030 249.400 ;
        RECT  30.440 247.660 64.400 249.400 ;
        RECT  0.600 124.090 64.400 129.850 ;
        RECT  1.640 124.090 63.600 135.790 ;
        RECT  1.810 124.090 2.830 154.520 ;
        RECT  4.040 123.970 60.900 171.560 ;
        RECT  1.640 155.040 63.600 171.560 ;
        RECT  1.640 183.580 63.600 185.950 ;
        RECT  5.490 124.090 63.600 200.820 ;
        RECT  1.640 196.170 63.600 200.820 ;
        RECT  56.930 123.970 57.210 201.060 ;
        RECT  0.600 0.600 64.400 60.480 ;
        RECT  2.000 0.000 63.000 88.700 ;
        RECT  0.600 0.600 1.480 91.220 ;
        RECT  0.600 90.750 64.400 91.220 ;
        LAYER TOP_M ;
        RECT  0.600 247.690 64.400 248.850 ;
        RECT  0.600 247.690 24.140 249.400 ;
        RECT  27.600 247.690 28.140 249.400 ;
        RECT  30.330 247.690 64.400 249.400 ;
        RECT  2.000 0.000 63.000 91.190 ;
        RECT  0.600 0.600 64.400 91.190 ;
    END
END pc3d01

MACRO pc3d00
    CLASS PAD ;
    FOREIGN pc3d00 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 65.000 BY 250.000 ;
    SYMMETRY X Y R90 ;
    SITE IOSite_c ;
    PIN PAD
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 55.440  LAYER TOP_M  ;
        ANTENNAPARTIALMETALSIDEAREA 294.161  LAYER M3  ;
        ANTENNAPARTIALMETALSIDEAREA 480.740  LAYER M2  ;
        ANTENNADIFFAREA 2657.280  LAYER TOP_M  ;
        ANTENNADIFFAREA 2657.280  LAYER M3  ;
        ANTENNADIFFAREA 1209.600  LAYER M2  ;
        ANTENNAPARTIALCUTAREA 632.318  LAYER TOP_V  ;
        ANTENNAPARTIALCUTAREA 349.898  LAYER V3  ;
        ANTENNAPARTIALCUTAREA 255.798  LAYER V2  ;
        PORT
        LAYER M3 ;
        RECT  21.430 247.650 31.230 250.000 ;
        LAYER M2 ;
        RECT  2.000 61.000 63.000 90.230 ;
        RECT  21.430 245.900 31.230 250.000 ;
        END
    END PAD
    PIN PADR
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 67.310  LAYER M1  ;
        ANTENNAPARTIALMETALSIDEAREA 35.658  LAYER M3  ;
        ANTENNAPARTIALMETALSIDEAREA 109.721  LAYER M2  ;
        ANTENNADIFFAREA 184.200  LAYER M3  ;
        ANTENNAPARTIALCUTAREA 0.338  LAYER V2  ;
        ANTENNAPARTIALCUTAREA 0.135  LAYER V3  ;
        PORT
        LAYER M3 ;
        RECT  33.230 249.270 34.310 250.000 ;
        LAYER M2 ;
        RECT  33.230 249.270 34.310 250.000 ;
        END
    END PADR
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        PORT
        LAYER M3 ;
        RECT  64.200 130.690 65.000 148.880 ;
        RECT  0.000 130.690 0.800 148.880 ;
        LAYER TOP_M ;
        RECT  0.000 123.850 65.000 154.560 ;
        LAYER M2 ;
        RECT  0.000 136.310 65.000 146.340 ;
        END
    END VSS
    PIN VSSO
        DIRECTION INOUT ;
        USE ground ;
        PORT
        LAYER M3 ;
        RECT  0.000 92.060 65.000 123.250 ;
        RECT  64.200 149.940 65.000 162.610 ;
        RECT  0.000 149.940 0.800 162.610 ;
        LAYER TOP_M ;
        RECT  0.000 92.060 65.000 123.250 ;
        RECT  0.000 155.410 65.000 162.610 ;
        LAYER M2 ;
        RECT  0.000 147.040 65.000 154.520 ;
        END
    END VSSO
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        PORT
        LAYER M3 ;
        RECT  64.200 163.510 65.000 190.890 ;
        RECT  0.000 163.510 0.800 190.890 ;
        LAYER TOP_M ;
        RECT  0.000 163.500 65.000 194.560 ;
        LAYER M2 ;
        RECT  0.000 172.080 65.000 183.060 ;
        END
    END VDD
    PIN VDDO
        DIRECTION INOUT ;
        USE power ;
        PORT
        LAYER M3 ;
        RECT  64.200 192.330 65.000 200.640 ;
        RECT  0.000 201.660 65.000 221.520 ;
        RECT  0.000 222.720 65.000 246.820 ;
        RECT  0.000 192.330 0.800 200.640 ;
        LAYER TOP_M ;
        RECT  0.000 195.170 65.000 200.640 ;
        RECT  0.000 201.660 65.000 221.520 ;
        RECT  0.000 222.720 65.000 246.820 ;
        LAYER M2 ;
        RECT  0.000 186.470 65.000 195.650 ;
        END
    END VDDO
    OBS
        LAYER M1 ;
        RECT  2.000 0.000 63.000 250.000 ;
        RECT  0.000 88.990 65.000 130.360 ;
        RECT  0.000 136.510 65.000 157.550 ;
        RECT  0.300 158.930 64.700 159.230 ;
        RECT  0.300 159.530 64.700 159.830 ;
        RECT  0.300 160.130 64.700 160.430 ;
        RECT  0.300 160.730 64.700 161.030 ;
        RECT  0.300 161.330 64.700 161.630 ;
        RECT  0.300 161.910 64.700 162.190 ;
        RECT  0.300 162.490 64.700 162.770 ;
        RECT  0.300 163.070 64.700 163.350 ;
        RECT  0.300 163.650 64.700 163.950 ;
        RECT  0.300 164.250 64.700 164.550 ;
        RECT  0.300 164.850 64.700 165.150 ;
        RECT  0.300 165.450 64.700 165.750 ;
        RECT  0.300 166.050 64.700 166.350 ;
        RECT  0.300 166.650 64.700 166.960 ;
        RECT  0.300 167.260 64.700 167.560 ;
        RECT  0.300 167.860 64.700 168.160 ;
        RECT  0.000 169.150 65.000 197.240 ;
        RECT  0.600 0.600 64.400 250.000 ;
        RECT  0.000 198.470 65.000 250.000 ;
        LAYER M2 ;
        RECT  63.180 196.430 63.670 249.400 ;
        RECT  0.600 196.440 64.400 245.110 ;
        RECT  32.020 196.440 64.400 248.480 ;
        RECT  0.600 196.440 20.640 249.400 ;
        RECT  32.020 196.440 32.440 249.400 ;
        RECT  35.100 196.440 64.400 249.400 ;
        RECT  0.600 183.850 64.400 185.680 ;
        RECT  7.125 183.850 46.210 185.855 ;
        RECT  1.620 154.990 2.550 171.435 ;
        RECT  58.960 155.200 59.270 171.290 ;
        RECT  60.005 155.235 60.315 171.290 ;
        RECT  0.600 155.310 64.400 171.290 ;
        RECT  55.705 155.310 56.505 171.405 ;
        RECT  1.620 155.310 17.700 171.435 ;
        RECT  2.000 0.000 63.000 60.210 ;
        RECT  0.600 0.600 64.400 60.210 ;
        RECT  0.600 0.600 1.210 135.520 ;
        RECT  0.600 91.020 64.400 135.520 ;
        RECT  4.140 91.020 61.000 135.690 ;
        LAYER M3 ;
        RECT  0.600 247.660 20.590 249.400 ;
        RECT  32.070 247.660 64.400 248.430 ;
        RECT  32.070 247.660 32.390 249.400 ;
        RECT  35.150 247.660 64.400 249.400 ;
        RECT  0.600 124.090 64.400 129.850 ;
        RECT  1.640 124.090 63.600 135.790 ;
        RECT  1.810 124.090 2.830 154.520 ;
        RECT  3.810 124.070 61.040 171.560 ;
        RECT  1.640 155.040 63.600 171.560 ;
        RECT  4.075 124.070 61.040 185.950 ;
        RECT  1.640 183.580 63.600 185.950 ;
        RECT  5.340 124.090 63.600 200.820 ;
        RECT  1.640 196.170 63.600 200.820 ;
        RECT  0.600 0.600 64.400 60.480 ;
        RECT  2.000 0.000 63.000 88.700 ;
        RECT  0.600 0.600 1.480 91.220 ;
        RECT  0.600 90.750 64.400 91.220 ;
        LAYER TOP_M ;
        RECT  0.600 247.690 20.700 249.400 ;
        RECT  31.960 247.690 64.400 248.540 ;
        RECT  31.960 247.690 32.500 249.400 ;
        RECT  35.040 247.690 64.400 249.400 ;
        RECT  2.000 0.000 63.000 91.190 ;
        RECT  0.600 0.600 64.400 91.190 ;
    END
END pc3d00

MACRO pc3c04
    CLASS PAD ;
    FOREIGN pc3c04 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 65.000 BY 250.000 ;
    SYMMETRY X Y R90 ;
    SITE IOSite_c ;
    PIN CCLK
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 54.897  LAYER M2  ;
        ANTENNAPARTIALMETALSIDEAREA 38.096  LAYER M3  ;
        ANTENNADIFFAREA 0.462  LAYER M3  ;
        ANTENNAPARTIALCUTAREA 0.135  LAYER V3  ;
        ANTENNAGATEAREA 192.960  LAYER M3  ;
        PORT
        LAYER M3 ;
        RECT  13.210 249.110 13.870 250.000 ;
        LAYER M2 ;
        RECT  13.210 249.110 13.870 250.000 ;
        END
    END CCLK
    PIN CP
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 1160.181  LAYER M3  ;
        ANTENNADIFFAREA 739.840  LAYER M3  ;
        PORT
        LAYER M3 ;
        RECT  18.100 249.150 46.900 250.000 ;
        LAYER M2 ;
        RECT  14.470 249.110 50.890 250.000 ;
        END
    END CP
    PIN VDDO
        DIRECTION INOUT ;
        USE power ;
        PORT
        LAYER M3 ;
        RECT  64.200 199.630 65.000 200.640 ;
        RECT  64.370 192.330 65.000 200.640 ;
        RECT  0.000 201.660 65.000 221.520 ;
        RECT  0.000 222.720 65.000 246.820 ;
        RECT  0.000 192.330 0.800 200.640 ;
        LAYER M2 ;
        RECT  0.000 186.470 65.000 195.650 ;
        LAYER TOP_M ;
        RECT  0.000 195.170 65.000 200.640 ;
        RECT  0.000 201.660 65.000 221.520 ;
        RECT  0.000 222.720 65.000 246.820 ;
        END
    END VDDO
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        PORT
        LAYER M3 ;
        RECT  64.370 163.510 65.000 190.890 ;
        RECT  0.000 163.510 0.800 190.890 ;
        LAYER M2 ;
        RECT  0.000 172.080 65.000 183.060 ;
        LAYER TOP_M ;
        RECT  0.000 163.500 65.000 194.560 ;
        END
    END VDD
    PIN VSSO
        DIRECTION INOUT ;
        USE ground ;
        PORT
        LAYER M3 ;
        RECT  0.000 92.060 65.000 123.250 ;
        RECT  64.370 149.940 65.000 162.610 ;
        RECT  0.000 149.940 0.800 162.610 ;
        LAYER M2 ;
        RECT  0.000 147.040 65.000 154.520 ;
        LAYER TOP_M ;
        RECT  0.000 92.060 65.000 123.250 ;
        RECT  0.000 155.410 65.000 162.610 ;
        END
    END VSSO
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        PORT
        LAYER M3 ;
        RECT  64.370 130.690 65.000 148.880 ;
        RECT  0.000 130.690 0.800 148.880 ;
        LAYER M2 ;
        RECT  0.000 136.310 65.000 146.340 ;
        LAYER TOP_M ;
        RECT  0.000 123.850 65.000 154.560 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.000 88.990 65.000 130.360 ;
        RECT  0.000 136.510 65.000 157.550 ;
        RECT  0.600 0.600 64.400 250.000 ;
        RECT  0.000 198.470 65.000 250.000 ;
        LAYER M2 ;
        RECT  0.600 196.440 64.400 248.320 ;
        RECT  0.600 196.440 12.420 249.400 ;
        RECT  51.680 196.440 64.400 249.400 ;
        RECT  0.600 183.850 64.400 185.680 ;
        RECT  15.630 155.120 16.520 171.290 ;
        RECT  20.350 155.120 21.240 171.290 ;
        RECT  25.070 155.120 25.960 171.290 ;
        RECT  29.790 155.120 30.680 171.290 ;
        RECT  34.510 155.120 35.400 171.290 ;
        RECT  39.230 155.120 40.120 171.290 ;
        RECT  43.950 155.120 44.840 171.290 ;
        RECT  48.670 155.120 49.560 171.290 ;
        RECT  0.600 155.310 64.400 171.290 ;
        RECT  0.600 0.600 64.400 135.520 ;
        LAYER M3 ;
        RECT  0.600 247.660 64.400 248.270 ;
        RECT  14.710 247.660 64.400 248.310 ;
        RECT  14.710 247.660 17.260 248.590 ;
        RECT  47.740 247.660 64.400 248.590 ;
        RECT  0.600 247.660 12.370 249.400 ;
        RECT  51.410 247.660 64.400 249.400 ;
        RECT  0.600 124.090 64.400 129.850 ;
        RECT  1.640 124.090 63.530 135.790 ;
        RECT  1.850 124.090 4.230 154.570 ;
        RECT  6.700 124.090 50.360 200.820 ;
        RECT  1.640 155.040 63.530 171.560 ;
        RECT  52.200 136.570 57.260 200.820 ;
        RECT  6.700 155.040 57.260 200.820 ;
        RECT  1.640 183.580 63.530 185.950 ;
        RECT  6.700 183.580 62.500 200.820 ;
        RECT  1.640 196.170 63.530 198.790 ;
        RECT  1.640 196.170 63.360 200.820 ;
        RECT  59.400 155.040 62.500 201.030 ;
        RECT  0.600 0.600 64.400 91.220 ;
        LAYER TOP_M ;
        RECT  0.600 247.690 64.400 248.380 ;
        RECT  14.600 247.690 64.400 248.420 ;
        RECT  0.600 247.690 12.480 249.400 ;
        RECT  14.600 247.690 17.370 249.400 ;
        RECT  47.630 247.690 64.400 249.400 ;
        RECT  0.600 0.600 64.400 91.190 ;
    END
END pc3c04

MACRO pc3c03
    CLASS PAD ;
    FOREIGN pc3c03 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 65.000 BY 250.000 ;
    SYMMETRY X Y R90 ;
    SITE IOSite_c ;
    PIN CP
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 760.815  LAYER M3  ;
        ANTENNADIFFAREA 369.920  LAYER M3  ;
        PORT
        LAYER M3 ;
        RECT  18.100 249.150 46.900 250.000 ;
        LAYER M2 ;
        RECT  14.470 247.680 50.890 250.000 ;
        RECT  42.150 198.490 50.890 250.000 ;
        RECT  32.950 208.740 50.890 250.000 ;
        RECT  14.470 208.740 32.050 250.000 ;
        RECT  14.470 198.430 22.850 250.000 ;
        END
    END CP
    PIN CCLK
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 54.897  LAYER M2  ;
        ANTENNAPARTIALMETALSIDEAREA 38.096  LAYER M3  ;
        ANTENNADIFFAREA 0.462  LAYER M3  ;
        ANTENNAPARTIALCUTAREA 0.135  LAYER V3  ;
        ANTENNAGATEAREA 96.480  LAYER M3  ;
        PORT
        LAYER M3 ;
        RECT  13.210 249.110 13.870 250.000 ;
        LAYER M2 ;
        RECT  13.210 249.110 13.870 250.000 ;
        END
    END CCLK
    PIN VDDO
        DIRECTION INOUT ;
        USE power ;
        PORT
        LAYER M3 ;
        RECT  64.200 199.630 65.000 200.640 ;
        RECT  64.370 192.330 65.000 200.640 ;
        RECT  0.000 201.660 65.000 221.520 ;
        RECT  0.000 222.720 65.000 246.820 ;
        RECT  0.000 192.330 0.800 200.640 ;
        LAYER M2 ;
        RECT  0.000 186.470 65.000 195.650 ;
        LAYER TOP_M ;
        RECT  0.000 195.170 65.000 200.640 ;
        RECT  0.000 201.660 65.000 221.520 ;
        RECT  0.000 222.720 65.000 246.820 ;
        END
    END VDDO
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        PORT
        LAYER M3 ;
        RECT  64.370 163.510 65.000 190.890 ;
        RECT  0.000 163.510 0.800 190.890 ;
        LAYER M2 ;
        RECT  0.000 172.080 65.000 183.060 ;
        LAYER TOP_M ;
        RECT  0.000 163.500 65.000 194.560 ;
        END
    END VDD
    PIN VSSO
        DIRECTION INOUT ;
        USE ground ;
        PORT
        LAYER M3 ;
        RECT  0.000 92.060 65.000 123.250 ;
        RECT  64.370 149.940 65.000 162.610 ;
        RECT  0.000 149.940 0.800 162.610 ;
        LAYER M2 ;
        RECT  0.000 147.040 65.000 154.520 ;
        LAYER TOP_M ;
        RECT  0.000 92.060 65.000 123.250 ;
        RECT  0.000 155.410 65.000 162.610 ;
        END
    END VSSO
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        PORT
        LAYER M3 ;
        RECT  64.370 130.690 65.000 148.880 ;
        RECT  0.000 130.690 0.800 148.880 ;
        LAYER M2 ;
        RECT  0.000 136.310 65.000 146.340 ;
        LAYER TOP_M ;
        RECT  0.000 123.850 65.000 154.560 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.000 88.990 65.000 130.360 ;
        RECT  0.000 136.510 65.000 157.550 ;
        RECT  0.600 0.600 64.400 250.000 ;
        RECT  0.000 198.470 65.000 250.000 ;
        LAYER M2 ;
        RECT  0.600 196.440 64.400 197.640 ;
        RECT  23.640 196.440 64.400 197.700 ;
        RECT  23.640 196.440 41.360 207.950 ;
        RECT  24.700 196.440 26.160 208.140 ;
        RECT  29.420 196.440 30.880 208.140 ;
        RECT  34.140 196.440 35.600 208.140 ;
        RECT  38.860 196.440 40.320 208.140 ;
        RECT  0.600 196.440 13.870 248.320 ;
        RECT  0.600 196.440 12.420 249.400 ;
        RECT  51.680 196.440 64.400 249.400 ;
        RECT  0.600 183.850 64.400 185.680 ;
        RECT  25.070 155.120 25.960 171.290 ;
        RECT  29.790 155.120 30.680 171.290 ;
        RECT  34.510 155.120 35.400 171.290 ;
        RECT  39.230 155.120 40.120 171.290 ;
        RECT  0.600 155.310 64.400 171.290 ;
        RECT  0.600 0.600 64.400 135.520 ;
        LAYER M3 ;
        RECT  0.600 247.660 13.950 248.270 ;
        RECT  0.600 247.660 12.370 249.400 ;
        RECT  51.410 247.660 64.400 249.400 ;
        RECT  0.600 124.090 64.400 129.850 ;
        RECT  1.640 124.090 63.530 135.790 ;
        RECT  1.850 124.090 4.230 154.570 ;
        RECT  52.200 136.570 57.260 200.820 ;
        RECT  1.640 155.040 63.530 171.560 ;
        RECT  1.640 183.580 63.530 185.950 ;
        RECT  6.700 183.580 62.500 197.910 ;
        RECT  6.700 124.090 50.890 197.910 ;
        RECT  23.370 155.040 57.260 197.970 ;
        RECT  51.410 196.170 63.530 198.790 ;
        RECT  14.470 124.090 22.850 200.070 ;
        RECT  42.150 124.090 50.890 200.070 ;
        RECT  1.640 196.170 13.950 200.820 ;
        RECT  23.370 124.090 41.630 200.820 ;
        RECT  51.410 196.170 63.360 200.820 ;
        RECT  59.400 155.040 62.500 201.030 ;
        RECT  0.600 0.600 64.400 91.220 ;
        LAYER TOP_M ;
        RECT  0.600 247.690 64.400 248.380 ;
        RECT  14.600 247.690 64.400 248.420 ;
        RECT  0.600 247.690 12.480 249.400 ;
        RECT  14.600 247.690 17.370 249.400 ;
        RECT  47.630 247.690 64.400 249.400 ;
        RECT  0.600 0.600 64.400 91.190 ;
    END
END pc3c03

MACRO pc3c02
    CLASS PAD ;
    FOREIGN pc3c02 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 65.000 BY 250.000 ;
    SYMMETRY X Y R90 ;
    SITE IOSite_c ;
    PIN CP
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 488.183  LAYER M3  ;
        ANTENNADIFFAREA 184.960  LAYER M3  ;
        PORT
        LAYER M3 ;
        RECT  18.100 249.150 46.900 250.000 ;
        LAYER M2 ;
        RECT  14.470 247.680 50.890 250.000 ;
        RECT  42.150 198.490 50.890 250.000 ;
        RECT  32.950 208.740 50.890 250.000 ;
        RECT  14.470 208.740 32.050 250.000 ;
        RECT  14.470 198.430 22.850 250.000 ;
        END
    END CP
    PIN CCLK
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 54.897  LAYER M2  ;
        ANTENNAPARTIALMETALSIDEAREA 38.096  LAYER M3  ;
        ANTENNADIFFAREA 0.462  LAYER M3  ;
        ANTENNAPARTIALCUTAREA 0.135  LAYER V3  ;
        ANTENNAGATEAREA 48.240  LAYER M3  ;
        PORT
        LAYER M3 ;
        RECT  13.210 249.110 13.870 250.000 ;
        LAYER M2 ;
        RECT  13.210 249.110 13.870 250.000 ;
        END
    END CCLK
    PIN VDDO
        DIRECTION INOUT ;
        USE power ;
        PORT
        LAYER M3 ;
        RECT  64.200 199.630 65.000 200.640 ;
        RECT  64.370 192.330 65.000 200.640 ;
        RECT  0.000 201.660 65.000 221.520 ;
        RECT  0.000 222.720 65.000 246.820 ;
        RECT  0.000 192.330 0.800 200.640 ;
        LAYER M2 ;
        RECT  0.000 186.470 65.000 195.650 ;
        LAYER TOP_M ;
        RECT  0.000 195.170 65.000 200.640 ;
        RECT  0.000 201.660 65.000 221.520 ;
        RECT  0.000 222.720 65.000 246.820 ;
        END
    END VDDO
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        PORT
        LAYER M3 ;
        RECT  64.370 163.510 65.000 190.890 ;
        RECT  0.000 163.510 0.800 190.890 ;
        LAYER M2 ;
        RECT  0.000 172.080 65.000 183.060 ;
        LAYER TOP_M ;
        RECT  0.000 163.500 65.000 194.560 ;
        END
    END VDD
    PIN VSSO
        DIRECTION INOUT ;
        USE ground ;
        PORT
        LAYER M3 ;
        RECT  0.000 92.060 65.000 123.250 ;
        RECT  64.370 149.940 65.000 162.610 ;
        RECT  0.000 149.940 0.800 162.610 ;
        LAYER M2 ;
        RECT  0.000 147.040 65.000 154.520 ;
        LAYER TOP_M ;
        RECT  0.000 92.060 65.000 123.250 ;
        RECT  0.000 155.410 65.000 162.610 ;
        END
    END VSSO
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        PORT
        LAYER M3 ;
        RECT  64.370 130.690 65.000 148.880 ;
        RECT  0.000 130.690 0.800 148.880 ;
        LAYER M2 ;
        RECT  0.000 136.310 65.000 146.340 ;
        LAYER TOP_M ;
        RECT  0.000 123.850 65.000 154.560 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.000 88.990 65.000 130.360 ;
        RECT  0.000 136.510 65.000 157.550 ;
        RECT  0.600 0.600 64.400 250.000 ;
        RECT  0.000 198.470 65.000 250.000 ;
        LAYER M2 ;
        RECT  0.600 196.440 64.400 197.640 ;
        RECT  23.640 196.440 64.400 197.700 ;
        RECT  23.640 196.440 41.360 207.950 ;
        RECT  29.420 196.440 30.880 208.140 ;
        RECT  34.140 196.440 35.600 208.140 ;
        RECT  0.600 196.440 13.870 248.320 ;
        RECT  0.600 196.440 12.420 249.400 ;
        RECT  51.680 196.440 64.400 249.400 ;
        RECT  0.600 183.850 64.400 185.680 ;
        RECT  29.790 155.120 30.680 171.290 ;
        RECT  34.510 155.120 35.400 171.290 ;
        RECT  0.600 155.310 64.400 171.290 ;
        RECT  0.600 0.600 64.400 135.520 ;
        LAYER M3 ;
        RECT  0.600 247.660 13.950 248.270 ;
        RECT  0.600 247.660 12.370 249.400 ;
        RECT  51.410 247.660 64.400 249.400 ;
        RECT  0.600 124.090 64.400 129.850 ;
        RECT  1.640 124.090 63.530 135.790 ;
        RECT  1.850 124.090 4.230 154.570 ;
        RECT  52.200 136.570 57.260 200.820 ;
        RECT  1.640 155.040 63.530 171.560 ;
        RECT  1.640 183.580 63.530 185.950 ;
        RECT  6.700 183.580 62.500 197.910 ;
        RECT  6.700 124.090 50.890 197.910 ;
        RECT  14.470 155.040 57.260 197.970 ;
        RECT  51.410 196.170 63.530 198.790 ;
        RECT  14.470 124.090 50.890 200.070 ;
        RECT  1.640 196.170 13.950 200.820 ;
        RECT  23.370 124.090 41.630 200.820 ;
        RECT  51.410 196.170 63.360 200.820 ;
        RECT  59.400 155.040 62.500 201.030 ;
        RECT  0.600 0.600 64.400 91.220 ;
        LAYER TOP_M ;
        RECT  0.600 247.690 64.400 248.380 ;
        RECT  14.600 247.690 64.400 248.420 ;
        RECT  0.600 247.690 12.480 249.400 ;
        RECT  14.600 247.690 17.370 249.400 ;
        RECT  47.630 247.690 64.400 249.400 ;
        RECT  0.600 0.600 64.400 91.190 ;
    END
END pc3c02

MACRO pc3c01
    CLASS PAD ;
    FOREIGN pc3c01 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 65.000 BY 250.000 ;
    SYMMETRY X Y R90 ;
    SITE IOSite_c ;
    PIN CP
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 352.630  LAYER M3  ;
        ANTENNADIFFAREA 92.480  LAYER M3  ;
        PORT
        LAYER M3 ;
        RECT  18.100 249.150 46.900 250.000 ;
        LAYER M2 ;
        RECT  14.470 249.110 50.890 250.000 ;
        END
    END CP
    PIN CCLK
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 54.897  LAYER M2  ;
        ANTENNAPARTIALMETALSIDEAREA 38.096  LAYER M3  ;
        ANTENNADIFFAREA 0.462  LAYER M3  ;
        ANTENNAPARTIALCUTAREA 0.135  LAYER V3  ;
        ANTENNAGATEAREA 24.120  LAYER M3  ;
        PORT
        LAYER M3 ;
        RECT  13.210 249.110 13.870 250.000 ;
        LAYER M2 ;
        RECT  13.210 249.110 13.870 250.000 ;
        END
    END CCLK
    PIN VDDO
        DIRECTION INOUT ;
        USE power ;
        PORT
        LAYER M3 ;
        RECT  64.200 199.630 65.000 200.640 ;
        RECT  64.370 192.330 65.000 200.640 ;
        RECT  0.000 201.660 65.000 221.520 ;
        RECT  0.000 222.720 65.000 246.820 ;
        RECT  0.000 192.330 0.800 200.640 ;
        LAYER M2 ;
        RECT  0.000 186.470 65.000 195.650 ;
        LAYER TOP_M ;
        RECT  0.000 195.170 65.000 200.640 ;
        RECT  0.000 201.660 65.000 221.520 ;
        RECT  0.000 222.720 65.000 246.820 ;
        END
    END VDDO
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        PORT
        LAYER M3 ;
        RECT  64.370 163.510 65.000 190.890 ;
        RECT  0.000 163.510 0.800 190.890 ;
        LAYER M2 ;
        RECT  0.000 172.080 65.000 183.060 ;
        LAYER TOP_M ;
        RECT  0.000 163.500 65.000 194.560 ;
        END
    END VDD
    PIN VSSO
        DIRECTION INOUT ;
        USE ground ;
        PORT
        LAYER M3 ;
        RECT  0.000 92.060 65.000 123.250 ;
        RECT  64.370 149.940 65.000 162.610 ;
        RECT  0.000 149.940 0.800 162.610 ;
        LAYER M2 ;
        RECT  0.000 147.040 65.000 154.520 ;
        LAYER TOP_M ;
        RECT  0.000 92.060 65.000 123.250 ;
        RECT  0.000 155.410 65.000 162.610 ;
        END
    END VSSO
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        PORT
        LAYER M3 ;
        RECT  64.370 130.690 65.000 148.880 ;
        RECT  0.000 130.690 0.800 148.880 ;
        LAYER M2 ;
        RECT  0.000 136.310 65.000 146.340 ;
        LAYER TOP_M ;
        RECT  0.000 123.850 65.000 154.560 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  0.000 88.990 65.000 130.360 ;
        RECT  0.000 136.510 65.000 157.550 ;
        RECT  0.600 0.600 64.400 250.000 ;
        RECT  0.000 198.470 65.000 250.000 ;
        LAYER M2 ;
        RECT  0.600 196.440 64.400 248.320 ;
        RECT  0.600 196.440 12.420 249.400 ;
        RECT  51.680 196.440 64.400 249.400 ;
        RECT  0.600 183.850 64.400 185.680 ;
        RECT  32.150 155.120 33.040 171.290 ;
        RECT  0.600 155.310 64.400 171.290 ;
        RECT  0.600 0.600 64.400 135.520 ;
        LAYER M3 ;
        RECT  0.600 247.660 64.400 248.270 ;
        RECT  14.710 247.660 64.400 248.310 ;
        RECT  14.710 247.660 17.260 248.590 ;
        RECT  47.740 247.660 64.400 248.590 ;
        RECT  0.600 247.660 12.370 249.400 ;
        RECT  51.410 247.660 64.400 249.400 ;
        RECT  0.600 124.090 64.400 129.850 ;
        RECT  1.640 124.090 63.530 135.790 ;
        RECT  1.850 124.090 4.230 154.570 ;
        RECT  6.700 124.090 50.890 200.820 ;
        RECT  1.640 155.040 63.530 171.560 ;
        RECT  52.200 136.570 57.260 200.820 ;
        RECT  6.700 155.040 57.260 200.820 ;
        RECT  1.640 183.580 63.530 185.950 ;
        RECT  6.700 183.580 62.500 200.820 ;
        RECT  1.640 196.170 63.530 198.790 ;
        RECT  1.640 196.170 63.360 200.820 ;
        RECT  59.400 155.040 62.500 201.030 ;
        RECT  0.600 0.600 64.400 91.220 ;
        LAYER TOP_M ;
        RECT  0.600 247.690 64.400 248.380 ;
        RECT  14.600 247.690 64.400 248.420 ;
        RECT  0.600 247.690 12.480 249.400 ;
        RECT  14.600 247.690 17.370 249.400 ;
        RECT  47.630 247.690 64.400 249.400 ;
        RECT  0.600 0.600 64.400 91.190 ;
    END
END pc3c01

MACRO pc3b25eu
    CLASS PAD ;
    FOREIGN pc3b25eu 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 65.000 BY 250.000 ;
    SYMMETRY X Y R90 ;
    SITE IOSite_c ;
    PIN PAD
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 55.440  LAYER TOP_M  ;
        ANTENNAPARTIALMETALSIDEAREA 287.938  LAYER M3  ;
        ANTENNAPARTIALMETALSIDEAREA 480.740  LAYER M2  ;
        ANTENNADIFFAREA 2657.280  LAYER TOP_M  ;
        ANTENNADIFFAREA 2657.280  LAYER M3  ;
        ANTENNADIFFAREA 1209.600  LAYER M2  ;
        ANTENNAPARTIALCUTAREA 632.318  LAYER TOP_V  ;
        ANTENNAPARTIALCUTAREA 349.898  LAYER V3  ;
        ANTENNAPARTIALCUTAREA 255.798  LAYER V2  ;
        PORT
        LAYER M3 ;
        RECT  23.740 249.580 25.740 250.000 ;
        LAYER M2 ;
        RECT  2.000 61.000 63.000 90.230 ;
        RECT  23.740 246.275 25.740 250.000 ;
        END
    END PAD
    PIN RENB
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 82.012  LAYER M2  ;
        ANTENNAPARTIALMETALSIDEAREA 44.266  LAYER M3  ;
        ANTENNADIFFAREA 1.000  LAYER M3  ;
        ANTENNAPARTIALCUTAREA 0.135  LAYER V3  ;
        ANTENNAGATEAREA 6.316  LAYER M3  ;
        PORT
        LAYER M3 ;
        RECT  30.930 249.580 31.660 250.000 ;
        LAYER M2 ;
        RECT  30.930 249.580 31.660 250.000 ;
        END
    END RENB
    PIN OEN
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 67.480  LAYER M3  ;
        ANTENNAPARTIALMETALSIDEAREA 67.374  LAYER M1  ;
        ANTENNAPARTIALMETALSIDEAREA 79.336  LAYER M2  ;
        ANTENNADIFFAREA 0.250  LAYER M3  ;
        ANTENNAPARTIALCUTAREA 0.135  LAYER V3  ;
        ANTENNAPARTIALCUTAREA 0.338  LAYER V2  ;
        ANTENNAGATEAREA 9.900  LAYER M3  ;
        ANTENNAGATEAREA 8.100  LAYER M2  ;
        PORT
        LAYER M3 ;
        RECT  29.900 249.580 30.630 250.000 ;
        LAYER M2 ;
        RECT  29.900 249.580 30.630 250.000 ;
        END
    END OEN
    PIN CIN
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 40.964  LAYER M3  ;
        ANTENNAPARTIALMETALSIDEAREA 67.374  LAYER M1  ;
        ANTENNAPARTIALMETALSIDEAREA 79.134  LAYER M2  ;
        ANTENNADIFFAREA 21.470  LAYER M3  ;
        ANTENNAPARTIALCUTAREA 0.203  LAYER V2  ;
        ANTENNAPARTIALCUTAREA 0.135  LAYER V3  ;
        PORT
        LAYER M3 ;
        RECT  28.870 249.580 29.600 250.000 ;
        LAYER M2 ;
        RECT  28.870 249.580 29.600 250.000 ;
        END
    END CIN
    PIN I
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 67.374  LAYER M1  ;
        ANTENNAPARTIALMETALSIDEAREA 79.415  LAYER M2  ;
        ANTENNAPARTIALMETALSIDEAREA 42.050  LAYER M3  ;
        ANTENNADIFFAREA 0.250  LAYER M3  ;
        ANTENNAPARTIALCUTAREA 0.270  LAYER V2  ;
        ANTENNAPARTIALCUTAREA 0.135  LAYER V3  ;
        ANTENNAGATEAREA 18.900  LAYER M2  ;
        ANTENNAGATEAREA 20.700  LAYER M3  ;
        PORT
        LAYER M3 ;
        RECT  27.840 249.580 28.570 250.000 ;
        LAYER M2 ;
        RECT  27.840 249.580 28.570 250.000 ;
        END
    END I
    PIN VDDO
        DIRECTION INOUT ;
        USE power ;
        PORT
        LAYER M3 ;
        RECT  64.200 192.330 65.000 200.640 ;
        RECT  0.000 201.660 65.000 221.520 ;
        RECT  0.000 222.720 65.000 246.820 ;
        RECT  0.000 192.330 0.800 200.640 ;
        LAYER M2 ;
        RECT  0.000 186.470 65.000 195.650 ;
        LAYER TOP_M ;
        RECT  0.000 195.170 65.000 200.640 ;
        RECT  0.000 201.660 65.000 221.520 ;
        RECT  0.000 222.720 65.000 246.820 ;
        END
    END VDDO
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        PORT
        LAYER M3 ;
        RECT  64.200 163.510 65.000 190.890 ;
        RECT  0.000 163.510 0.800 190.890 ;
        LAYER M2 ;
        RECT  0.000 172.080 65.000 183.060 ;
        LAYER TOP_M ;
        RECT  0.000 163.500 65.000 194.560 ;
        END
    END VDD
    PIN VSSO
        DIRECTION INOUT ;
        USE ground ;
        PORT
        LAYER M3 ;
        RECT  0.000 92.060 65.000 123.250 ;
        RECT  64.200 149.940 65.000 162.610 ;
        RECT  0.000 149.940 0.800 162.610 ;
        LAYER M2 ;
        RECT  0.000 147.040 65.000 154.520 ;
        LAYER TOP_M ;
        RECT  0.000 92.060 65.000 123.250 ;
        RECT  0.000 155.410 65.000 162.610 ;
        END
    END VSSO
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        PORT
        LAYER M3 ;
        RECT  64.200 130.690 65.000 148.880 ;
        RECT  0.000 130.690 0.800 148.880 ;
        LAYER M2 ;
        RECT  0.000 136.310 65.000 146.340 ;
        LAYER TOP_M ;
        RECT  0.000 123.850 65.000 154.560 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  2.000 0.000 63.000 250.000 ;
        RECT  0.000 88.990 65.000 130.360 ;
        RECT  0.000 136.510 65.000 157.550 ;
        RECT  0.300 158.330 64.700 158.630 ;
        RECT  0.300 158.930 64.700 159.230 ;
        RECT  0.300 159.530 64.700 159.830 ;
        RECT  0.300 160.130 64.700 160.430 ;
        RECT  0.300 160.730 64.700 161.030 ;
        RECT  0.300 161.330 64.700 161.630 ;
        RECT  0.300 161.910 64.700 162.190 ;
        RECT  0.300 162.490 64.700 162.770 ;
        RECT  0.300 163.070 64.700 163.350 ;
        RECT  0.300 163.650 64.700 163.950 ;
        RECT  0.300 164.250 64.700 164.550 ;
        RECT  0.300 164.850 64.700 165.150 ;
        RECT  0.300 165.450 64.700 165.750 ;
        RECT  0.300 166.050 64.700 166.350 ;
        RECT  0.300 166.650 64.700 166.960 ;
        RECT  0.300 167.260 64.700 167.560 ;
        RECT  0.300 167.860 64.700 168.160 ;
        RECT  0.000 169.150 65.000 197.240 ;
        RECT  0.600 0.600 64.400 250.000 ;
        RECT  0.000 198.470 65.000 250.000 ;
        LAYER M2 ;
        RECT  1.740 196.420 2.020 249.400 ;
        RECT  63.180 196.430 63.670 249.400 ;
        RECT  0.600 196.440 64.400 245.485 ;
        RECT  26.530 196.440 64.400 248.790 ;
        RECT  0.600 196.440 22.950 249.400 ;
        RECT  26.530 196.440 27.050 249.400 ;
        RECT  32.450 196.440 64.400 249.400 ;
        RECT  18.260 183.720 52.060 185.680 ;
        RECT  55.990 183.710 56.310 185.880 ;
        RECT  0.600 183.850 64.400 185.680 ;
        RECT  46.230 183.720 51.730 185.870 ;
        RECT  53.850 183.850 54.840 185.870 ;
        RECT  55.375 183.850 61.350 185.880 ;
        RECT  4.480 154.920 7.530 171.290 ;
        RECT  8.170 155.125 8.490 171.290 ;
        RECT  20.200 155.160 20.550 171.290 ;
        RECT  20.830 155.140 21.150 171.290 ;
        RECT  22.525 155.200 22.815 171.290 ;
        RECT  24.440 155.120 24.720 171.290 ;
        RECT  25.000 155.240 25.280 171.290 ;
        RECT  32.590 155.120 36.460 171.290 ;
        RECT  48.830 155.120 49.150 171.290 ;
        RECT  49.530 155.120 49.810 171.290 ;
        RECT  50.115 155.125 50.445 171.290 ;
        RECT  51.780 155.120 53.325 171.290 ;
        RECT  53.690 155.110 53.990 171.325 ;
        RECT  57.750 155.130 58.030 171.290 ;
        RECT  0.600 155.310 64.400 171.290 ;
        RECT  23.850 155.310 24.130 171.310 ;
        RECT  53.050 155.310 57.845 171.325 ;
        RECT  23.290 155.310 23.570 171.330 ;
        RECT  46.995 155.310 47.380 171.375 ;
        RECT  3.170 155.310 3.450 171.380 ;
        RECT  33.350 155.310 39.255 171.480 ;
        RECT  41.100 155.310 43.485 171.480 ;
        RECT  60.160 155.310 63.000 171.480 ;
        RECT  2.000 0.000 63.000 60.210 ;
        RECT  0.600 0.600 64.400 60.210 ;
        RECT  0.600 0.600 1.210 135.520 ;
        RECT  0.600 91.020 64.400 135.520 ;
        RECT  4.080 91.020 60.940 135.690 ;
        RECT  62.580 91.020 62.995 135.710 ;
        LAYER M3 ;
        RECT  0.600 247.660 23.220 248.740 ;
        RECT  0.600 247.660 22.900 249.400 ;
        RECT  26.260 247.660 64.400 248.740 ;
        RECT  26.580 247.660 27.000 249.400 ;
        RECT  32.500 247.660 64.400 249.400 ;
        RECT  4.040 123.970 60.900 200.820 ;
        RECT  0.600 124.090 64.400 129.850 ;
        RECT  1.640 124.090 63.600 135.790 ;
        RECT  1.810 124.090 2.830 154.520 ;
        RECT  1.640 155.040 63.600 171.560 ;
        RECT  1.640 183.580 63.600 185.950 ;
        RECT  2.860 155.040 63.600 200.820 ;
        RECT  3.510 124.090 63.600 200.820 ;
        RECT  1.640 196.170 63.600 200.820 ;
        RECT  54.265 123.970 54.545 201.060 ;
        RECT  0.600 0.600 64.400 60.480 ;
        RECT  2.000 0.000 63.000 88.700 ;
        RECT  0.600 0.600 1.480 91.220 ;
        RECT  0.600 90.750 64.400 91.220 ;
        LAYER TOP_M ;
        RECT  0.600 247.690 64.400 248.850 ;
        RECT  0.600 247.690 23.010 249.400 ;
        RECT  26.470 247.690 27.110 249.400 ;
        RECT  32.390 247.690 64.400 249.400 ;
        RECT  2.000 0.000 63.000 91.190 ;
        RECT  0.600 0.600 64.400 91.190 ;
    END
END pc3b25eu

MACRO pc3b21eu
    CLASS PAD ;
    FOREIGN pc3b21eu 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 65.000 BY 250.000 ;
    SYMMETRY X Y R90 ;
    SITE IOSite_c ;
    PIN RENB
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 82.012  LAYER M2  ;
        ANTENNAPARTIALMETALSIDEAREA 44.266  LAYER M3  ;
        ANTENNADIFFAREA 1.000  LAYER M3  ;
        ANTENNAPARTIALCUTAREA 0.135  LAYER V3  ;
        ANTENNAGATEAREA 6.316  LAYER M3  ;
        PORT
        LAYER M3 ;
        RECT  30.930 249.580 31.660 250.000 ;
        LAYER M2 ;
        RECT  30.930 249.580 31.660 250.000 ;
        END
    END RENB
    PIN PAD
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 55.440  LAYER TOP_M  ;
        ANTENNAPARTIALMETALSIDEAREA 287.938  LAYER M3  ;
        ANTENNAPARTIALMETALSIDEAREA 480.740  LAYER M2  ;
        ANTENNADIFFAREA 2657.280  LAYER TOP_M  ;
        ANTENNADIFFAREA 2657.280  LAYER M3  ;
        ANTENNADIFFAREA 1209.600  LAYER M2  ;
        ANTENNAPARTIALCUTAREA 632.318  LAYER TOP_V  ;
        ANTENNAPARTIALCUTAREA 349.898  LAYER V3  ;
        ANTENNAPARTIALCUTAREA 255.798  LAYER V2  ;
        PORT
        LAYER M3 ;
        RECT  23.740 249.580 25.740 250.000 ;
        LAYER M2 ;
        RECT  2.000 61.000 63.000 90.230 ;
        RECT  23.740 246.275 25.740 250.000 ;
        END
    END PAD
    PIN CIN
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 79.134  LAYER M2  ;
        ANTENNAPARTIALMETALSIDEAREA 67.374  LAYER M1  ;
        ANTENNAPARTIALMETALSIDEAREA 40.964  LAYER M3  ;
        ANTENNADIFFAREA 21.470  LAYER M3  ;
        ANTENNAPARTIALCUTAREA 0.135  LAYER V3  ;
        ANTENNAPARTIALCUTAREA 0.203  LAYER V2  ;
        PORT
        LAYER M3 ;
        RECT  28.870 249.580 29.600 250.000 ;
        LAYER M2 ;
        RECT  28.870 249.580 29.600 250.000 ;
        END
    END CIN
    PIN OEN
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 79.336  LAYER M2  ;
        ANTENNAPARTIALMETALSIDEAREA 67.374  LAYER M1  ;
        ANTENNAPARTIALMETALSIDEAREA 67.480  LAYER M3  ;
        ANTENNADIFFAREA 0.250  LAYER M3  ;
        ANTENNAPARTIALCUTAREA 0.338  LAYER V2  ;
        ANTENNAPARTIALCUTAREA 0.135  LAYER V3  ;
        ANTENNAGATEAREA 8.100  LAYER M2  ;
        ANTENNAGATEAREA 9.900  LAYER M3  ;
        PORT
        LAYER M3 ;
        RECT  29.900 249.580 30.630 250.000 ;
        LAYER M2 ;
        RECT  29.900 249.580 30.630 250.000 ;
        END
    END OEN
    PIN I
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 67.374  LAYER M1  ;
        ANTENNAPARTIALMETALSIDEAREA 79.415  LAYER M2  ;
        ANTENNAPARTIALMETALSIDEAREA 42.050  LAYER M3  ;
        ANTENNADIFFAREA 0.250  LAYER M3  ;
        ANTENNAPARTIALCUTAREA 0.203  LAYER V2  ;
        ANTENNAPARTIALCUTAREA 0.135  LAYER V3  ;
        ANTENNAGATEAREA 8.100  LAYER M2  ;
        ANTENNAGATEAREA 9.900  LAYER M3  ;
        PORT
        LAYER M3 ;
        RECT  27.840 249.580 28.570 250.000 ;
        LAYER M2 ;
        RECT  27.840 249.580 28.570 250.000 ;
        END
    END I
    PIN VDDO
        DIRECTION INOUT ;
        USE power ;
        PORT
        LAYER M3 ;
        RECT  64.200 192.330 65.000 200.640 ;
        RECT  0.000 201.660 65.000 221.520 ;
        RECT  0.000 222.720 65.000 246.820 ;
        RECT  0.000 192.330 0.800 200.640 ;
        LAYER M2 ;
        RECT  0.000 186.470 65.000 195.650 ;
        LAYER TOP_M ;
        RECT  0.000 195.170 65.000 200.640 ;
        RECT  0.000 201.660 65.000 221.520 ;
        RECT  0.000 222.720 65.000 246.820 ;
        END
    END VDDO
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        PORT
        LAYER M3 ;
        RECT  64.200 163.510 65.000 190.890 ;
        RECT  0.000 163.510 0.800 190.890 ;
        LAYER M2 ;
        RECT  0.000 172.080 65.000 183.060 ;
        LAYER TOP_M ;
        RECT  0.000 163.500 65.000 194.560 ;
        END
    END VDD
    PIN VSSO
        DIRECTION INOUT ;
        USE ground ;
        PORT
        LAYER M3 ;
        RECT  0.000 92.060 65.000 123.250 ;
        RECT  64.200 149.940 65.000 162.610 ;
        RECT  0.000 149.940 0.800 162.610 ;
        LAYER M2 ;
        RECT  0.000 147.040 65.000 154.520 ;
        LAYER TOP_M ;
        RECT  0.000 92.060 65.000 123.250 ;
        RECT  0.000 155.410 65.000 162.610 ;
        END
    END VSSO
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        PORT
        LAYER M3 ;
        RECT  64.200 130.690 65.000 148.880 ;
        RECT  0.000 130.690 0.800 148.880 ;
        LAYER M2 ;
        RECT  0.000 136.310 65.000 146.340 ;
        LAYER TOP_M ;
        RECT  0.000 123.850 65.000 154.560 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  2.000 0.000 63.000 250.000 ;
        RECT  0.000 88.990 65.000 130.360 ;
        RECT  0.000 136.510 65.000 157.550 ;
        RECT  0.300 158.330 64.700 158.630 ;
        RECT  0.300 158.930 64.700 159.230 ;
        RECT  0.300 159.530 64.700 159.830 ;
        RECT  0.300 160.130 64.700 160.430 ;
        RECT  0.300 160.730 64.700 161.030 ;
        RECT  0.300 161.330 64.700 161.630 ;
        RECT  0.300 161.910 64.700 162.190 ;
        RECT  0.300 162.490 64.700 162.770 ;
        RECT  0.300 163.070 64.700 163.350 ;
        RECT  0.300 163.650 64.700 163.950 ;
        RECT  0.300 164.250 64.700 164.550 ;
        RECT  0.300 164.850 64.700 165.150 ;
        RECT  0.300 165.450 64.700 165.750 ;
        RECT  0.300 166.050 64.700 166.350 ;
        RECT  0.300 166.650 64.700 166.960 ;
        RECT  0.300 167.260 64.700 167.560 ;
        RECT  0.300 167.860 64.700 168.160 ;
        RECT  0.000 169.150 65.000 197.240 ;
        RECT  0.600 0.600 64.400 250.000 ;
        RECT  0.000 198.470 65.000 250.000 ;
        LAYER M2 ;
        RECT  1.740 196.420 2.020 249.400 ;
        RECT  63.180 196.430 63.670 249.400 ;
        RECT  0.600 196.440 64.400 245.485 ;
        RECT  26.530 196.440 64.400 248.790 ;
        RECT  0.600 196.440 22.950 249.400 ;
        RECT  26.530 196.440 27.050 249.400 ;
        RECT  32.450 196.440 64.400 249.400 ;
        RECT  17.025 183.720 52.380 185.680 ;
        RECT  55.995 183.710 56.315 185.880 ;
        RECT  0.600 183.850 64.400 185.680 ;
        RECT  46.230 183.720 51.730 185.870 ;
        RECT  53.850 183.850 54.840 185.870 ;
        RECT  55.375 183.850 61.350 185.880 ;
        RECT  19.375 155.200 19.665 171.290 ;
        RECT  21.290 155.120 21.570 171.290 ;
        RECT  21.850 155.240 22.130 171.290 ;
        RECT  22.410 155.160 22.760 171.290 ;
        RECT  23.060 155.140 23.380 171.290 ;
        RECT  48.835 155.120 49.155 171.290 ;
        RECT  49.535 155.120 49.815 171.290 ;
        RECT  50.120 155.125 50.450 171.290 ;
        RECT  51.785 155.120 53.330 171.290 ;
        RECT  53.695 155.110 53.995 171.325 ;
        RECT  57.755 155.130 58.035 171.290 ;
        RECT  0.600 155.310 64.400 171.290 ;
        RECT  20.700 155.310 20.980 171.310 ;
        RECT  53.055 155.310 57.850 171.325 ;
        RECT  20.140 155.310 20.420 171.330 ;
        RECT  46.850 155.310 47.235 171.375 ;
        RECT  3.220 155.310 3.500 171.380 ;
        RECT  33.970 155.310 39.260 171.480 ;
        RECT  41.105 155.310 43.490 171.480 ;
        RECT  60.015 155.310 62.855 171.480 ;
        RECT  2.000 0.000 63.000 60.210 ;
        RECT  0.600 0.600 64.400 60.210 ;
        RECT  0.600 0.600 1.210 135.520 ;
        RECT  0.600 91.020 64.400 135.520 ;
        RECT  4.080 91.020 60.940 135.690 ;
        RECT  62.580 91.020 62.995 135.710 ;
        LAYER M3 ;
        RECT  0.600 247.660 23.220 248.740 ;
        RECT  0.600 247.660 22.900 249.400 ;
        RECT  26.260 247.660 64.400 248.740 ;
        RECT  26.580 247.660 27.000 249.400 ;
        RECT  32.500 247.660 64.400 249.400 ;
        RECT  0.600 124.090 64.400 129.850 ;
        RECT  3.990 123.970 60.900 135.790 ;
        RECT  1.640 124.090 63.600 135.790 ;
        RECT  1.810 124.090 2.830 154.520 ;
        RECT  1.640 155.040 63.600 171.560 ;
        RECT  1.640 183.580 63.600 185.950 ;
        RECT  2.910 155.040 63.600 200.820 ;
        RECT  5.155 124.090 63.600 200.820 ;
        RECT  1.640 196.170 63.600 200.820 ;
        RECT  54.265 123.970 54.545 201.060 ;
        RECT  0.600 0.600 64.400 60.480 ;
        RECT  2.000 0.000 63.000 88.700 ;
        RECT  0.600 0.600 1.480 91.220 ;
        RECT  0.600 90.750 64.400 91.220 ;
        LAYER TOP_M ;
        RECT  0.600 247.690 64.400 248.850 ;
        RECT  0.600 247.690 23.010 249.400 ;
        RECT  26.470 247.690 27.110 249.400 ;
        RECT  32.390 247.690 64.400 249.400 ;
        RECT  2.000 0.000 63.000 91.190 ;
        RECT  0.600 0.600 64.400 91.190 ;
    END
END pc3b21eu

MACRO pc3b05u
    CLASS PAD ;
    FOREIGN pc3b05u 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 65.000 BY 250.000 ;
    SYMMETRY X Y R90 ;
    SITE IOSite_c ;
    PIN PAD
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 55.440  LAYER TOP_M  ;
        ANTENNAPARTIALMETALSIDEAREA 287.938  LAYER M3  ;
        ANTENNAPARTIALMETALSIDEAREA 480.740  LAYER M2  ;
        ANTENNADIFFAREA 2657.280  LAYER TOP_M  ;
        ANTENNADIFFAREA 2657.280  LAYER M3  ;
        ANTENNADIFFAREA 1209.600  LAYER M2  ;
        ANTENNAPARTIALCUTAREA 632.318  LAYER TOP_V  ;
        ANTENNAPARTIALCUTAREA 349.898  LAYER V3  ;
        ANTENNAPARTIALCUTAREA 255.798  LAYER V2  ;
        PORT
        LAYER M3 ;
        RECT  23.740 249.580 25.740 250.000 ;
        LAYER M2 ;
        RECT  2.000 61.000 63.000 90.230 ;
        RECT  23.740 246.275 25.740 250.000 ;
        END
    END PAD
    PIN CIN
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 32.277  LAYER M3  ;
        ANTENNAPARTIALMETALSIDEAREA 96.916  LAYER M2  ;
        ANTENNAPARTIALMETALSIDEAREA 67.374  LAYER M1  ;
        ANTENNADIFFAREA 20.600  LAYER M3  ;
        ANTENNAPARTIALCUTAREA 0.135  LAYER V3  ;
        ANTENNAPARTIALCUTAREA 0.203  LAYER V2  ;
        PORT
        LAYER M3 ;
        RECT  28.870 249.580 29.600 250.000 ;
        LAYER M2 ;
        RECT  28.870 249.580 29.600 250.000 ;
        END
    END CIN
    PIN OEN
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 80.634  LAYER M2  ;
        ANTENNAPARTIALMETALSIDEAREA 67.374  LAYER M1  ;
        ANTENNAPARTIALMETALSIDEAREA 41.679  LAYER M3  ;
        ANTENNADIFFAREA 0.250  LAYER M3  ;
        ANTENNAPARTIALCUTAREA 0.203  LAYER V2  ;
        ANTENNAPARTIALCUTAREA 0.135  LAYER V3  ;
        ANTENNAGATEAREA 8.100  LAYER M2  ;
        ANTENNAGATEAREA 9.900  LAYER M3  ;
        PORT
        LAYER M3 ;
        RECT  29.900 249.580 30.630 250.000 ;
        LAYER M2 ;
        RECT  29.900 249.580 30.630 250.000 ;
        END
    END OEN
    PIN I
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 67.374  LAYER M1  ;
        ANTENNAPARTIALMETALSIDEAREA 80.804  LAYER M2  ;
        ANTENNAPARTIALMETALSIDEAREA 41.096  LAYER M3  ;
        ANTENNADIFFAREA 0.250  LAYER M3  ;
        ANTENNAPARTIALCUTAREA 0.270  LAYER V2  ;
        ANTENNAPARTIALCUTAREA 0.135  LAYER V3  ;
        ANTENNAGATEAREA 18.900  LAYER M2  ;
        ANTENNAGATEAREA 20.700  LAYER M3  ;
        PORT
        LAYER M3 ;
        RECT  27.840 249.580 28.570 250.000 ;
        LAYER M2 ;
        RECT  27.840 249.580 28.570 250.000 ;
        END
    END I
    PIN VDDO
        DIRECTION INOUT ;
        USE power ;
        PORT
        LAYER M3 ;
        RECT  64.200 192.330 65.000 200.640 ;
        RECT  0.000 201.660 65.000 221.520 ;
        RECT  0.000 222.720 65.000 246.820 ;
        RECT  0.000 192.330 0.800 200.640 ;
        LAYER M2 ;
        RECT  0.000 186.470 65.000 195.650 ;
        LAYER TOP_M ;
        RECT  0.000 195.170 65.000 200.640 ;
        RECT  0.000 201.660 65.000 221.520 ;
        RECT  0.000 222.720 65.000 246.820 ;
        END
    END VDDO
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        PORT
        LAYER M3 ;
        RECT  64.200 163.510 65.000 190.890 ;
        RECT  0.000 163.510 0.800 190.890 ;
        LAYER M2 ;
        RECT  0.000 172.080 65.000 183.060 ;
        LAYER TOP_M ;
        RECT  0.000 163.500 65.000 194.560 ;
        END
    END VDD
    PIN VSSO
        DIRECTION INOUT ;
        USE ground ;
        PORT
        LAYER M3 ;
        RECT  0.000 92.060 65.000 123.250 ;
        RECT  64.200 149.940 65.000 162.610 ;
        RECT  0.000 149.940 0.800 162.610 ;
        LAYER M2 ;
        RECT  0.000 147.040 65.000 154.520 ;
        LAYER TOP_M ;
        RECT  0.000 92.060 65.000 123.250 ;
        RECT  0.000 155.410 65.000 162.610 ;
        END
    END VSSO
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        PORT
        LAYER M3 ;
        RECT  64.200 130.690 65.000 148.880 ;
        RECT  0.000 130.690 0.800 148.880 ;
        LAYER M2 ;
        RECT  0.000 136.310 65.000 146.340 ;
        LAYER TOP_M ;
        RECT  0.000 123.850 65.000 154.560 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  2.000 0.000 63.000 250.000 ;
        RECT  0.000 88.990 65.000 130.360 ;
        RECT  0.000 136.510 65.000 157.550 ;
        RECT  0.315 158.150 64.700 158.460 ;
        RECT  0.300 158.930 64.700 159.230 ;
        RECT  0.300 159.530 64.700 159.830 ;
        RECT  0.300 160.130 64.700 160.430 ;
        RECT  0.300 160.730 64.700 161.030 ;
        RECT  0.300 161.330 64.700 161.630 ;
        RECT  0.300 161.910 64.700 162.190 ;
        RECT  0.300 162.490 64.700 162.770 ;
        RECT  0.300 163.070 64.700 163.350 ;
        RECT  0.300 163.650 64.700 163.950 ;
        RECT  0.300 164.250 64.700 164.550 ;
        RECT  0.300 164.850 64.700 165.150 ;
        RECT  0.300 165.450 64.700 165.750 ;
        RECT  0.300 166.050 64.700 166.350 ;
        RECT  0.300 166.650 64.700 166.960 ;
        RECT  0.300 167.260 64.700 167.560 ;
        RECT  0.300 167.860 64.700 168.160 ;
        RECT  0.000 169.150 65.000 197.240 ;
        RECT  0.600 0.600 64.400 250.000 ;
        RECT  0.000 198.470 65.000 250.000 ;
        LAYER M2 ;
        RECT  1.840 196.420 2.120 249.400 ;
        RECT  63.180 196.430 63.670 249.400 ;
        RECT  0.600 196.440 64.400 245.485 ;
        RECT  26.530 196.440 64.400 248.790 ;
        RECT  0.600 196.440 22.950 249.400 ;
        RECT  26.530 196.440 27.050 249.400 ;
        RECT  31.420 196.440 64.400 249.400 ;
        RECT  19.440 183.720 52.225 185.680 ;
        RECT  0.600 183.850 64.400 185.680 ;
        RECT  46.230 183.720 51.730 185.870 ;
        RECT  55.235 183.850 56.645 185.900 ;
        RECT  4.480 154.920 7.530 171.290 ;
        RECT  8.170 155.125 8.490 171.290 ;
        RECT  22.160 155.160 22.510 171.290 ;
        RECT  22.810 155.140 23.130 171.290 ;
        RECT  31.960 155.120 35.830 171.290 ;
        RECT  53.655 155.035 53.935 171.290 ;
        RECT  56.365 155.280 56.645 171.315 ;
        RECT  57.120 155.300 57.400 171.315 ;
        RECT  57.835 155.130 58.115 171.315 ;
        RECT  0.600 155.310 64.400 171.290 ;
        RECT  56.240 155.310 61.880 171.315 ;
        RECT  53.895 155.310 55.870 171.370 ;
        RECT  3.170 155.310 3.450 171.380 ;
        RECT  34.655 155.310 38.715 171.480 ;
        RECT  39.605 155.310 42.020 171.480 ;
        RECT  2.000 0.000 63.000 60.210 ;
        RECT  0.600 0.600 64.400 60.210 ;
        RECT  0.600 0.600 1.210 135.520 ;
        RECT  0.600 91.020 64.400 135.520 ;
        RECT  4.080 91.020 60.940 135.690 ;
        RECT  62.580 91.020 62.995 135.710 ;
        LAYER M3 ;
        RECT  0.600 247.660 23.220 248.740 ;
        RECT  0.600 247.660 22.900 249.400 ;
        RECT  26.260 247.660 64.400 248.740 ;
        RECT  26.580 247.660 27.000 249.400 ;
        RECT  31.470 247.660 64.400 249.400 ;
        RECT  0.600 124.090 64.400 129.850 ;
        RECT  1.640 124.090 63.600 135.790 ;
        RECT  1.810 124.090 2.830 154.520 ;
        RECT  3.510 124.090 63.600 171.560 ;
        RECT  4.040 123.970 60.900 171.560 ;
        RECT  1.640 155.040 63.600 171.560 ;
        RECT  1.640 183.580 63.600 185.950 ;
        RECT  5.515 124.090 63.600 200.820 ;
        RECT  1.640 196.170 63.600 200.820 ;
        RECT  56.300 123.970 56.580 201.060 ;
        RECT  0.600 0.600 64.400 60.480 ;
        RECT  2.000 0.000 63.000 88.700 ;
        RECT  0.600 0.600 1.480 91.220 ;
        RECT  0.600 90.750 64.400 91.220 ;
        LAYER TOP_M ;
        RECT  0.600 247.690 64.400 248.850 ;
        RECT  0.600 247.690 23.010 249.400 ;
        RECT  26.470 247.690 27.110 249.400 ;
        RECT  31.360 247.690 64.400 249.400 ;
        RECT  2.000 0.000 63.000 91.190 ;
        RECT  0.600 0.600 64.400 91.190 ;
    END
END pc3b05u

MACRO pc3b05d
    CLASS PAD ;
    FOREIGN pc3b05d 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 65.000 BY 250.000 ;
    SYMMETRY X Y R90 ;
    SITE IOSite_c ;
    PIN PAD
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 55.440  LAYER TOP_M  ;
        ANTENNAPARTIALMETALSIDEAREA 287.938  LAYER M3  ;
        ANTENNAPARTIALMETALSIDEAREA 480.740  LAYER M2  ;
        ANTENNADIFFAREA 2657.280  LAYER TOP_M  ;
        ANTENNADIFFAREA 2657.280  LAYER M3  ;
        ANTENNADIFFAREA 1209.600  LAYER M2  ;
        ANTENNAPARTIALCUTAREA 632.318  LAYER TOP_V  ;
        ANTENNAPARTIALCUTAREA 349.898  LAYER V3  ;
        ANTENNAPARTIALCUTAREA 255.798  LAYER V2  ;
        PORT
        LAYER M3 ;
        RECT  23.740 249.580 25.740 250.000 ;
        LAYER M2 ;
        RECT  2.000 61.000 63.000 90.230 ;
        RECT  23.740 246.275 25.740 250.000 ;
        END
    END PAD
    PIN CIN
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 32.277  LAYER M3  ;
        ANTENNAPARTIALMETALSIDEAREA 96.916  LAYER M2  ;
        ANTENNAPARTIALMETALSIDEAREA 67.374  LAYER M1  ;
        ANTENNADIFFAREA 20.600  LAYER M3  ;
        ANTENNAPARTIALCUTAREA 0.135  LAYER V3  ;
        ANTENNAPARTIALCUTAREA 0.203  LAYER V2  ;
        PORT
        LAYER M3 ;
        RECT  28.870 249.580 29.600 250.000 ;
        LAYER M2 ;
        RECT  28.870 249.580 29.600 250.000 ;
        END
    END CIN
    PIN OEN
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 80.634  LAYER M2  ;
        ANTENNAPARTIALMETALSIDEAREA 67.374  LAYER M1  ;
        ANTENNAPARTIALMETALSIDEAREA 41.679  LAYER M3  ;
        ANTENNADIFFAREA 0.250  LAYER M3  ;
        ANTENNAPARTIALCUTAREA 0.203  LAYER V2  ;
        ANTENNAPARTIALCUTAREA 0.135  LAYER V3  ;
        ANTENNAGATEAREA 8.100  LAYER M2  ;
        ANTENNAGATEAREA 9.900  LAYER M3  ;
        PORT
        LAYER M3 ;
        RECT  29.900 249.580 30.630 250.000 ;
        LAYER M2 ;
        RECT  29.900 249.580 30.630 250.000 ;
        END
    END OEN
    PIN I
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 67.374  LAYER M1  ;
        ANTENNAPARTIALMETALSIDEAREA 80.804  LAYER M2  ;
        ANTENNAPARTIALMETALSIDEAREA 41.096  LAYER M3  ;
        ANTENNADIFFAREA 0.250  LAYER M3  ;
        ANTENNAPARTIALCUTAREA 0.270  LAYER V2  ;
        ANTENNAPARTIALCUTAREA 0.135  LAYER V3  ;
        ANTENNAGATEAREA 18.900  LAYER M2  ;
        ANTENNAGATEAREA 20.700  LAYER M3  ;
        PORT
        LAYER M3 ;
        RECT  27.840 249.580 28.570 250.000 ;
        LAYER M2 ;
        RECT  27.840 249.580 28.570 250.000 ;
        END
    END I
    PIN VDDO
        DIRECTION INOUT ;
        USE power ;
        PORT
        LAYER M3 ;
        RECT  64.200 192.330 65.000 200.640 ;
        RECT  0.000 201.660 65.000 221.520 ;
        RECT  0.000 222.720 65.000 246.820 ;
        RECT  0.000 192.330 0.800 200.640 ;
        LAYER M2 ;
        RECT  0.000 186.470 65.000 195.650 ;
        LAYER TOP_M ;
        RECT  0.000 195.170 65.000 200.640 ;
        RECT  0.000 201.660 65.000 221.520 ;
        RECT  0.000 222.720 65.000 246.820 ;
        END
    END VDDO
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        PORT
        LAYER M3 ;
        RECT  64.200 163.510 65.000 190.890 ;
        RECT  0.000 163.510 0.800 190.890 ;
        LAYER M2 ;
        RECT  0.000 172.080 65.000 183.060 ;
        LAYER TOP_M ;
        RECT  0.000 163.500 65.000 194.560 ;
        END
    END VDD
    PIN VSSO
        DIRECTION INOUT ;
        USE ground ;
        PORT
        LAYER M3 ;
        RECT  0.000 92.060 65.000 123.250 ;
        RECT  64.200 149.940 65.000 162.610 ;
        RECT  0.000 149.940 0.800 162.610 ;
        LAYER M2 ;
        RECT  0.000 147.040 65.000 154.520 ;
        LAYER TOP_M ;
        RECT  0.000 92.060 65.000 123.250 ;
        RECT  0.000 155.410 65.000 162.610 ;
        END
    END VSSO
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        PORT
        LAYER M3 ;
        RECT  64.200 130.690 65.000 148.880 ;
        RECT  0.000 130.690 0.800 148.880 ;
        LAYER M2 ;
        RECT  0.000 136.310 65.000 146.340 ;
        LAYER TOP_M ;
        RECT  0.000 123.850 65.000 154.560 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  2.000 0.000 63.000 250.000 ;
        RECT  0.000 88.990 65.000 130.360 ;
        RECT  0.000 136.510 65.000 157.550 ;
        RECT  0.315 158.150 64.700 158.460 ;
        RECT  0.300 158.930 64.700 159.230 ;
        RECT  0.300 159.530 64.700 159.830 ;
        RECT  0.300 160.130 64.700 160.430 ;
        RECT  0.300 160.730 64.700 161.030 ;
        RECT  0.300 161.330 64.700 161.630 ;
        RECT  0.300 161.910 64.700 162.190 ;
        RECT  0.300 162.490 64.700 162.770 ;
        RECT  0.300 163.070 64.700 163.350 ;
        RECT  0.300 163.650 64.700 163.950 ;
        RECT  0.300 164.250 64.700 164.550 ;
        RECT  0.300 164.850 64.700 165.150 ;
        RECT  0.300 165.450 64.700 165.750 ;
        RECT  0.300 166.050 64.700 166.350 ;
        RECT  0.300 166.650 64.700 166.960 ;
        RECT  0.300 167.260 64.700 167.560 ;
        RECT  0.300 167.860 64.700 168.160 ;
        RECT  0.000 169.150 65.000 197.240 ;
        RECT  0.600 0.600 64.400 250.000 ;
        RECT  0.000 198.470 65.000 250.000 ;
        LAYER M2 ;
        RECT  1.840 196.420 2.120 249.400 ;
        RECT  63.180 196.430 63.670 249.400 ;
        RECT  0.600 196.440 64.400 245.485 ;
        RECT  26.530 196.440 64.400 248.790 ;
        RECT  0.600 196.440 22.950 249.400 ;
        RECT  26.530 196.440 27.050 249.400 ;
        RECT  31.420 196.440 64.400 249.400 ;
        RECT  19.440 183.720 52.225 185.680 ;
        RECT  0.600 183.850 64.400 185.680 ;
        RECT  46.230 183.720 51.730 185.870 ;
        RECT  55.235 183.850 56.645 185.900 ;
        RECT  4.480 154.920 7.530 171.290 ;
        RECT  8.170 155.125 8.490 171.290 ;
        RECT  22.160 155.160 22.510 171.290 ;
        RECT  22.810 155.140 23.130 171.290 ;
        RECT  31.960 155.120 35.830 171.290 ;
        RECT  49.195 155.130 51.435 171.290 ;
        RECT  52.375 155.300 52.685 171.290 ;
        RECT  53.655 155.035 53.935 171.290 ;
        RECT  56.365 155.280 56.645 171.315 ;
        RECT  57.120 155.300 57.400 171.315 ;
        RECT  57.835 155.130 58.115 171.315 ;
        RECT  0.600 155.310 64.400 171.290 ;
        RECT  56.240 155.310 61.880 171.315 ;
        RECT  53.895 155.310 55.870 171.370 ;
        RECT  3.170 155.310 3.450 171.380 ;
        RECT  34.655 155.310 38.715 171.480 ;
        RECT  39.605 155.310 42.020 171.480 ;
        RECT  2.000 0.000 63.000 60.210 ;
        RECT  0.600 0.600 64.400 60.210 ;
        RECT  0.600 0.600 1.210 135.520 ;
        RECT  0.600 91.020 64.400 135.520 ;
        RECT  4.080 91.020 60.940 135.690 ;
        RECT  62.580 91.020 62.995 135.710 ;
        LAYER M3 ;
        RECT  0.600 247.660 23.220 248.740 ;
        RECT  0.600 247.660 22.900 249.400 ;
        RECT  26.260 247.660 64.400 248.740 ;
        RECT  26.580 247.660 27.000 249.400 ;
        RECT  31.470 247.660 64.400 249.400 ;
        RECT  0.600 124.090 64.400 129.850 ;
        RECT  1.640 124.090 63.600 135.790 ;
        RECT  1.810 124.090 2.830 154.520 ;
        RECT  3.510 124.090 63.600 171.560 ;
        RECT  4.040 123.970 60.900 171.560 ;
        RECT  1.640 155.040 63.600 171.560 ;
        RECT  1.640 183.580 63.600 185.950 ;
        RECT  5.515 124.090 63.600 200.820 ;
        RECT  1.640 196.170 63.600 200.820 ;
        RECT  56.300 123.970 56.580 201.060 ;
        RECT  0.600 0.600 64.400 60.480 ;
        RECT  2.000 0.000 63.000 88.700 ;
        RECT  0.600 0.600 1.480 91.220 ;
        RECT  0.600 90.750 64.400 91.220 ;
        LAYER TOP_M ;
        RECT  0.600 247.690 64.400 248.850 ;
        RECT  0.600 247.690 23.010 249.400 ;
        RECT  26.470 247.690 27.110 249.400 ;
        RECT  31.360 247.690 64.400 249.400 ;
        RECT  2.000 0.000 63.000 91.190 ;
        RECT  0.600 0.600 64.400 91.190 ;
    END
END pc3b05d

MACRO pc3b05
    CLASS PAD ;
    FOREIGN pc3b05 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 65.000 BY 250.000 ;
    SYMMETRY X Y R90 ;
    SITE IOSite_c ;
    PIN PAD
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 55.440  LAYER TOP_M  ;
        ANTENNAPARTIALMETALSIDEAREA 287.938  LAYER M3  ;
        ANTENNAPARTIALMETALSIDEAREA 480.740  LAYER M2  ;
        ANTENNADIFFAREA 2657.280  LAYER TOP_M  ;
        ANTENNADIFFAREA 2657.280  LAYER M3  ;
        ANTENNADIFFAREA 1209.600  LAYER M2  ;
        ANTENNAPARTIALCUTAREA 632.318  LAYER TOP_V  ;
        ANTENNAPARTIALCUTAREA 349.898  LAYER V3  ;
        ANTENNAPARTIALCUTAREA 255.798  LAYER V2  ;
        PORT
        LAYER M3 ;
        RECT  23.740 249.580 25.740 250.000 ;
        LAYER M2 ;
        RECT  2.000 61.000 63.000 90.230 ;
        RECT  23.740 246.275 25.740 250.000 ;
        END
    END PAD
    PIN CIN
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 32.277  LAYER M3  ;
        ANTENNAPARTIALMETALSIDEAREA 96.916  LAYER M2  ;
        ANTENNAPARTIALMETALSIDEAREA 67.374  LAYER M1  ;
        ANTENNADIFFAREA 20.600  LAYER M3  ;
        ANTENNAPARTIALCUTAREA 0.135  LAYER V3  ;
        ANTENNAPARTIALCUTAREA 0.203  LAYER V2  ;
        PORT
        LAYER M3 ;
        RECT  28.870 249.580 29.600 250.000 ;
        LAYER M2 ;
        RECT  28.870 249.580 29.600 250.000 ;
        END
    END CIN
    PIN OEN
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 80.634  LAYER M2  ;
        ANTENNAPARTIALMETALSIDEAREA 67.374  LAYER M1  ;
        ANTENNAPARTIALMETALSIDEAREA 41.679  LAYER M3  ;
        ANTENNADIFFAREA 0.250  LAYER M3  ;
        ANTENNAPARTIALCUTAREA 0.203  LAYER V2  ;
        ANTENNAPARTIALCUTAREA 0.135  LAYER V3  ;
        ANTENNAGATEAREA 8.100  LAYER M2  ;
        ANTENNAGATEAREA 9.900  LAYER M3  ;
        PORT
        LAYER M3 ;
        RECT  29.900 249.580 30.630 250.000 ;
        LAYER M2 ;
        RECT  29.900 249.580 30.630 250.000 ;
        END
    END OEN
    PIN I
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 67.374  LAYER M1  ;
        ANTENNAPARTIALMETALSIDEAREA 80.804  LAYER M2  ;
        ANTENNAPARTIALMETALSIDEAREA 41.096  LAYER M3  ;
        ANTENNADIFFAREA 0.250  LAYER M3  ;
        ANTENNAPARTIALCUTAREA 0.270  LAYER V2  ;
        ANTENNAPARTIALCUTAREA 0.135  LAYER V3  ;
        ANTENNAGATEAREA 18.900  LAYER M2  ;
        ANTENNAGATEAREA 20.700  LAYER M3  ;
        PORT
        LAYER M3 ;
        RECT  27.840 249.580 28.570 250.000 ;
        LAYER M2 ;
        RECT  27.840 249.580 28.570 250.000 ;
        END
    END I
    PIN VDDO
        DIRECTION INOUT ;
        USE power ;
        PORT
        LAYER M3 ;
        RECT  64.200 192.330 65.000 200.640 ;
        RECT  0.000 201.660 65.000 221.520 ;
        RECT  0.000 222.720 65.000 246.820 ;
        RECT  0.000 192.330 0.800 200.640 ;
        LAYER M2 ;
        RECT  0.000 186.470 65.000 195.650 ;
        LAYER TOP_M ;
        RECT  0.000 195.170 65.000 200.640 ;
        RECT  0.000 201.660 65.000 221.520 ;
        RECT  0.000 222.720 65.000 246.820 ;
        END
    END VDDO
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        PORT
        LAYER M3 ;
        RECT  64.200 163.510 65.000 190.890 ;
        RECT  0.000 163.510 0.800 190.890 ;
        LAYER M2 ;
        RECT  0.000 172.080 65.000 183.060 ;
        LAYER TOP_M ;
        RECT  0.000 163.500 65.000 194.560 ;
        END
    END VDD
    PIN VSSO
        DIRECTION INOUT ;
        USE ground ;
        PORT
        LAYER M3 ;
        RECT  0.000 92.060 65.000 123.250 ;
        RECT  64.200 149.940 65.000 162.610 ;
        RECT  0.000 149.940 0.800 162.610 ;
        LAYER M2 ;
        RECT  0.000 147.040 65.000 154.520 ;
        LAYER TOP_M ;
        RECT  0.000 92.060 65.000 123.250 ;
        RECT  0.000 155.410 65.000 162.610 ;
        END
    END VSSO
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        PORT
        LAYER M3 ;
        RECT  64.200 130.690 65.000 148.880 ;
        RECT  0.000 130.690 0.800 148.880 ;
        LAYER M2 ;
        RECT  0.000 136.310 65.000 146.340 ;
        LAYER TOP_M ;
        RECT  0.000 123.850 65.000 154.560 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  2.000 0.000 63.000 250.000 ;
        RECT  0.000 88.990 65.000 130.360 ;
        RECT  0.000 136.510 65.000 157.550 ;
        RECT  0.315 158.150 64.700 158.460 ;
        RECT  0.300 158.930 64.700 159.230 ;
        RECT  0.300 159.530 64.700 159.830 ;
        RECT  0.300 160.130 64.700 160.430 ;
        RECT  0.300 160.730 64.700 161.030 ;
        RECT  0.300 161.330 64.700 161.630 ;
        RECT  0.300 161.910 64.700 162.190 ;
        RECT  0.300 162.490 64.700 162.770 ;
        RECT  0.300 163.070 64.700 163.350 ;
        RECT  0.300 163.650 64.700 163.950 ;
        RECT  0.300 164.250 64.700 164.550 ;
        RECT  0.300 164.850 64.700 165.150 ;
        RECT  0.300 165.450 64.700 165.750 ;
        RECT  0.300 166.050 64.700 166.350 ;
        RECT  0.300 166.650 64.700 166.960 ;
        RECT  0.300 167.260 64.700 167.560 ;
        RECT  0.300 167.860 64.700 168.160 ;
        RECT  0.000 169.150 65.000 197.240 ;
        RECT  0.600 0.600 64.400 250.000 ;
        RECT  0.000 198.470 65.000 250.000 ;
        LAYER M2 ;
        RECT  1.840 196.420 2.120 249.400 ;
        RECT  63.180 196.430 63.670 249.400 ;
        RECT  0.600 196.440 64.400 245.485 ;
        RECT  26.530 196.440 64.400 248.790 ;
        RECT  0.600 196.440 22.950 249.400 ;
        RECT  26.530 196.440 27.050 249.400 ;
        RECT  31.420 196.440 64.400 249.400 ;
        RECT  19.440 183.720 52.225 185.680 ;
        RECT  0.600 183.850 64.400 185.680 ;
        RECT  46.230 183.720 51.730 185.870 ;
        RECT  55.235 183.850 56.645 185.900 ;
        RECT  4.480 154.920 7.530 171.290 ;
        RECT  8.170 155.125 8.490 171.290 ;
        RECT  22.160 155.160 22.510 171.290 ;
        RECT  22.810 155.140 23.130 171.290 ;
        RECT  31.960 155.120 35.830 171.290 ;
        RECT  53.655 155.035 53.935 171.290 ;
        RECT  56.365 155.280 56.645 171.315 ;
        RECT  57.120 155.300 57.400 171.315 ;
        RECT  57.835 155.130 58.115 171.315 ;
        RECT  0.600 155.310 64.400 171.290 ;
        RECT  56.240 155.310 61.880 171.315 ;
        RECT  53.895 155.310 55.870 171.370 ;
        RECT  3.170 155.310 3.450 171.380 ;
        RECT  34.655 155.310 38.715 171.480 ;
        RECT  39.605 155.310 42.020 171.480 ;
        RECT  2.000 0.000 63.000 60.210 ;
        RECT  0.600 0.600 64.400 60.210 ;
        RECT  0.600 0.600 1.210 135.520 ;
        RECT  0.600 91.020 64.400 135.520 ;
        RECT  4.080 91.020 60.940 135.690 ;
        RECT  62.580 91.020 62.995 135.710 ;
        LAYER M3 ;
        RECT  0.600 247.660 23.220 248.740 ;
        RECT  0.600 247.660 22.900 249.400 ;
        RECT  26.260 247.660 64.400 248.740 ;
        RECT  26.580 247.660 27.000 249.400 ;
        RECT  31.470 247.660 64.400 249.400 ;
        RECT  0.600 124.090 64.400 129.850 ;
        RECT  1.640 124.090 63.600 135.790 ;
        RECT  1.810 124.090 2.830 154.520 ;
        RECT  3.510 124.090 63.600 171.560 ;
        RECT  4.040 123.970 60.900 171.560 ;
        RECT  1.640 155.040 63.600 171.560 ;
        RECT  1.640 183.580 63.600 185.950 ;
        RECT  5.515 124.090 63.600 200.820 ;
        RECT  1.640 196.170 63.600 200.820 ;
        RECT  56.300 123.970 56.580 201.060 ;
        RECT  0.600 0.600 64.400 60.480 ;
        RECT  2.000 0.000 63.000 88.700 ;
        RECT  0.600 0.600 1.480 91.220 ;
        RECT  0.600 90.750 64.400 91.220 ;
        LAYER TOP_M ;
        RECT  0.600 247.690 64.400 248.850 ;
        RECT  0.600 247.690 23.010 249.400 ;
        RECT  26.470 247.690 27.110 249.400 ;
        RECT  31.360 247.690 64.400 249.400 ;
        RECT  2.000 0.000 63.000 91.190 ;
        RECT  0.600 0.600 64.400 91.190 ;
    END
END pc3b05

MACRO pc3b04u
    CLASS PAD ;
    FOREIGN pc3b04u 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 65.000 BY 250.000 ;
    SYMMETRY X Y R90 ;
    SITE IOSite_c ;
    PIN PAD
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 55.440  LAYER TOP_M  ;
        ANTENNAPARTIALMETALSIDEAREA 287.938  LAYER M3  ;
        ANTENNAPARTIALMETALSIDEAREA 480.740  LAYER M2  ;
        ANTENNADIFFAREA 2657.280  LAYER TOP_M  ;
        ANTENNADIFFAREA 1209.600  LAYER M2  ;
        ANTENNADIFFAREA 2657.280  LAYER M3  ;
        ANTENNAPARTIALCUTAREA 632.318  LAYER TOP_V  ;
        ANTENNAPARTIALCUTAREA 349.898  LAYER V3  ;
        ANTENNAPARTIALCUTAREA 255.798  LAYER V2  ;
        PORT
        LAYER M3 ;
        RECT  23.740 249.580 25.740 250.000 ;
        LAYER M2 ;
        RECT  2.000 61.000 63.000 90.230 ;
        RECT  23.740 246.275 25.740 250.000 ;
        END
    END PAD
    PIN OEN
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 80.634  LAYER M2  ;
        ANTENNAPARTIALMETALSIDEAREA 41.679  LAYER M3  ;
        ANTENNAPARTIALMETALSIDEAREA 67.374  LAYER M1  ;
        ANTENNADIFFAREA 0.250  LAYER M3  ;
        ANTENNAPARTIALCUTAREA 0.203  LAYER V2  ;
        ANTENNAPARTIALCUTAREA 0.135  LAYER V3  ;
        ANTENNAGATEAREA 9.900  LAYER M3  ;
        ANTENNAGATEAREA 8.100  LAYER M2  ;
        PORT
        LAYER M3 ;
        RECT  29.900 249.580 30.630 250.000 ;
        LAYER M2 ;
        RECT  29.900 249.580 30.630 250.000 ;
        END
    END OEN
    PIN CIN
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 32.277  LAYER M3  ;
        ANTENNAPARTIALMETALSIDEAREA 96.916  LAYER M2  ;
        ANTENNAPARTIALMETALSIDEAREA 67.374  LAYER M1  ;
        ANTENNADIFFAREA 20.600  LAYER M3  ;
        ANTENNAPARTIALCUTAREA 0.135  LAYER V3  ;
        ANTENNAPARTIALCUTAREA 0.203  LAYER V2  ;
        PORT
        LAYER M3 ;
        RECT  28.870 249.580 29.600 250.000 ;
        LAYER M2 ;
        RECT  28.870 249.580 29.600 250.000 ;
        END
    END CIN
    PIN I
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 67.374  LAYER M1  ;
        ANTENNAPARTIALMETALSIDEAREA 80.804  LAYER M2  ;
        ANTENNAPARTIALMETALSIDEAREA 41.096  LAYER M3  ;
        ANTENNADIFFAREA 0.250  LAYER M3  ;
        ANTENNAPARTIALCUTAREA 0.270  LAYER V2  ;
        ANTENNAPARTIALCUTAREA 0.135  LAYER V3  ;
        ANTENNAGATEAREA 18.900  LAYER M2  ;
        ANTENNAGATEAREA 20.700  LAYER M3  ;
        PORT
        LAYER M3 ;
        RECT  27.840 249.580 28.570 250.000 ;
        LAYER M2 ;
        RECT  27.840 249.580 28.570 250.000 ;
        END
    END I
    PIN VSSO
        DIRECTION INOUT ;
        USE ground ;
        PORT
        LAYER M3 ;
        RECT  0.000 92.060 65.000 123.250 ;
        RECT  64.200 149.940 65.000 162.610 ;
        RECT  0.000 149.940 0.800 162.610 ;
        LAYER M2 ;
        RECT  0.000 147.040 65.000 154.520 ;
        LAYER TOP_M ;
        RECT  0.000 92.060 65.000 123.250 ;
        RECT  0.000 155.410 65.000 162.610 ;
        END
    END VSSO
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        PORT
        LAYER M3 ;
        RECT  64.200 130.690 65.000 148.880 ;
        RECT  0.000 130.690 0.800 148.880 ;
        LAYER M2 ;
        RECT  0.000 136.310 65.000 146.340 ;
        LAYER TOP_M ;
        RECT  0.000 123.850 65.000 154.560 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        PORT
        LAYER M3 ;
        RECT  64.200 163.510 65.000 190.890 ;
        RECT  0.000 163.510 0.800 190.890 ;
        LAYER M2 ;
        RECT  0.000 172.080 65.000 183.060 ;
        LAYER TOP_M ;
        RECT  0.000 163.500 65.000 194.560 ;
        END
    END VDD
    PIN VDDO
        DIRECTION INOUT ;
        USE power ;
        PORT
        LAYER M3 ;
        RECT  64.200 192.330 65.000 200.640 ;
        RECT  0.000 201.660 65.000 221.520 ;
        RECT  0.000 222.720 65.000 246.820 ;
        RECT  0.000 192.330 0.800 200.640 ;
        LAYER M2 ;
        RECT  0.000 186.470 65.000 195.650 ;
        LAYER TOP_M ;
        RECT  0.000 195.170 65.000 200.640 ;
        RECT  0.000 201.660 65.000 221.520 ;
        RECT  0.000 222.720 65.000 246.820 ;
        END
    END VDDO
    OBS
        LAYER M1 ;
        RECT  2.000 0.000 63.000 250.000 ;
        RECT  0.000 88.990 65.000 130.360 ;
        RECT  0.000 136.510 65.000 157.550 ;
        RECT  0.315 158.150 64.700 158.460 ;
        RECT  0.300 158.930 64.700 159.230 ;
        RECT  0.300 159.530 64.700 159.830 ;
        RECT  0.300 160.130 64.700 160.430 ;
        RECT  0.300 160.730 64.700 161.030 ;
        RECT  0.300 161.330 64.700 161.630 ;
        RECT  0.300 161.910 64.700 162.190 ;
        RECT  0.300 162.490 64.700 162.770 ;
        RECT  0.300 163.070 64.700 163.350 ;
        RECT  0.300 163.650 64.700 163.950 ;
        RECT  0.300 164.250 64.700 164.550 ;
        RECT  0.300 164.850 64.700 165.150 ;
        RECT  0.300 165.450 64.700 165.750 ;
        RECT  0.300 166.050 64.700 166.350 ;
        RECT  0.300 166.650 64.700 166.960 ;
        RECT  0.300 167.260 64.700 167.560 ;
        RECT  0.300 167.860 64.700 168.160 ;
        RECT  0.000 169.150 65.000 197.240 ;
        RECT  0.600 0.600 64.400 250.000 ;
        RECT  0.000 198.470 65.000 250.000 ;
        LAYER M2 ;
        RECT  1.840 196.420 2.120 249.400 ;
        RECT  63.180 196.430 63.670 249.400 ;
        RECT  0.600 196.440 64.400 245.485 ;
        RECT  26.530 196.440 64.400 248.790 ;
        RECT  0.600 196.440 22.950 249.400 ;
        RECT  26.530 196.440 27.050 249.400 ;
        RECT  31.420 196.440 64.400 249.400 ;
        RECT  19.140 183.720 52.180 185.680 ;
        RECT  0.600 183.850 64.400 185.680 ;
        RECT  55.195 183.850 56.950 185.850 ;
        RECT  46.230 183.720 51.730 185.870 ;
        RECT  4.830 155.120 7.380 171.290 ;
        RECT  8.170 155.125 8.490 171.290 ;
        RECT  22.160 155.160 22.510 171.290 ;
        RECT  22.810 155.140 23.130 171.290 ;
        RECT  53.655 155.035 53.935 171.290 ;
        RECT  56.365 155.280 56.645 171.315 ;
        RECT  57.120 155.300 57.400 171.315 ;
        RECT  57.835 155.130 58.115 171.315 ;
        RECT  0.600 155.310 64.400 171.290 ;
        RECT  56.240 155.310 61.880 171.315 ;
        RECT  53.895 155.310 55.870 171.370 ;
        RECT  33.575 155.310 34.075 171.375 ;
        RECT  3.175 155.310 3.455 171.380 ;
        RECT  34.655 155.310 38.715 171.480 ;
        RECT  39.605 155.310 42.020 171.480 ;
        RECT  2.000 0.000 63.000 60.210 ;
        RECT  0.600 0.600 64.400 60.210 ;
        RECT  0.600 0.600 1.210 135.520 ;
        RECT  0.600 91.020 64.400 135.520 ;
        RECT  4.080 91.020 60.940 135.690 ;
        RECT  62.580 91.020 62.995 135.710 ;
        LAYER M3 ;
        RECT  0.600 247.660 23.220 248.740 ;
        RECT  0.600 247.660 22.900 249.400 ;
        RECT  26.260 247.660 64.400 248.740 ;
        RECT  26.580 247.660 27.000 249.400 ;
        RECT  31.470 247.660 64.400 249.400 ;
        RECT  0.600 124.090 64.400 129.850 ;
        RECT  1.640 124.090 63.600 135.790 ;
        RECT  1.810 124.090 2.830 154.520 ;
        RECT  3.195 124.090 63.600 171.560 ;
        RECT  3.325 123.900 61.330 171.560 ;
        RECT  1.640 155.040 63.600 171.560 ;
        RECT  1.640 183.580 63.600 185.950 ;
        RECT  5.515 124.090 63.600 200.820 ;
        RECT  1.640 196.170 63.600 200.820 ;
        RECT  56.300 123.900 56.580 201.060 ;
        RECT  0.600 0.600 64.400 60.480 ;
        RECT  2.000 0.000 63.000 88.700 ;
        RECT  0.600 0.600 1.480 91.220 ;
        RECT  0.600 90.750 64.400 91.220 ;
        LAYER TOP_M ;
        RECT  0.600 247.690 64.400 248.850 ;
        RECT  0.600 247.690 23.010 249.400 ;
        RECT  26.470 247.690 27.110 249.400 ;
        RECT  31.360 247.690 64.400 249.400 ;
        RECT  2.000 0.000 63.000 91.190 ;
        RECT  0.600 0.600 64.400 91.190 ;
    END
END pc3b04u

MACRO pc3b04d
    CLASS PAD ;
    FOREIGN pc3b04d 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 65.000 BY 250.000 ;
    SYMMETRY X Y R90 ;
    SITE IOSite_c ;
    PIN PAD
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 55.440  LAYER TOP_M  ;
        ANTENNAPARTIALMETALSIDEAREA 287.938  LAYER M3  ;
        ANTENNAPARTIALMETALSIDEAREA 480.740  LAYER M2  ;
        ANTENNADIFFAREA 2657.280  LAYER TOP_M  ;
        ANTENNADIFFAREA 1209.600  LAYER M2  ;
        ANTENNADIFFAREA 2657.280  LAYER M3  ;
        ANTENNAPARTIALCUTAREA 632.318  LAYER TOP_V  ;
        ANTENNAPARTIALCUTAREA 349.898  LAYER V3  ;
        ANTENNAPARTIALCUTAREA 255.798  LAYER V2  ;
        PORT
        LAYER M3 ;
        RECT  23.740 249.580 25.740 250.000 ;
        LAYER M2 ;
        RECT  2.000 61.000 63.000 90.230 ;
        RECT  23.740 246.275 25.740 250.000 ;
        END
    END PAD
    PIN OEN
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 80.634  LAYER M2  ;
        ANTENNAPARTIALMETALSIDEAREA 41.679  LAYER M3  ;
        ANTENNAPARTIALMETALSIDEAREA 67.374  LAYER M1  ;
        ANTENNADIFFAREA 0.250  LAYER M3  ;
        ANTENNAPARTIALCUTAREA 0.203  LAYER V2  ;
        ANTENNAPARTIALCUTAREA 0.135  LAYER V3  ;
        ANTENNAGATEAREA 9.900  LAYER M3  ;
        ANTENNAGATEAREA 8.100  LAYER M2  ;
        PORT
        LAYER M3 ;
        RECT  29.900 249.580 30.630 250.000 ;
        LAYER M2 ;
        RECT  29.900 249.580 30.630 250.000 ;
        END
    END OEN
    PIN CIN
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 32.277  LAYER M3  ;
        ANTENNAPARTIALMETALSIDEAREA 96.916  LAYER M2  ;
        ANTENNAPARTIALMETALSIDEAREA 67.374  LAYER M1  ;
        ANTENNADIFFAREA 20.600  LAYER M3  ;
        ANTENNAPARTIALCUTAREA 0.135  LAYER V3  ;
        ANTENNAPARTIALCUTAREA 0.203  LAYER V2  ;
        PORT
        LAYER M3 ;
        RECT  28.870 249.580 29.600 250.000 ;
        LAYER M2 ;
        RECT  28.870 249.580 29.600 250.000 ;
        END
    END CIN
    PIN I
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 67.374  LAYER M1  ;
        ANTENNAPARTIALMETALSIDEAREA 80.804  LAYER M2  ;
        ANTENNAPARTIALMETALSIDEAREA 41.096  LAYER M3  ;
        ANTENNADIFFAREA 0.250  LAYER M3  ;
        ANTENNAPARTIALCUTAREA 0.270  LAYER V2  ;
        ANTENNAPARTIALCUTAREA 0.135  LAYER V3  ;
        ANTENNAGATEAREA 18.900  LAYER M2  ;
        ANTENNAGATEAREA 20.700  LAYER M3  ;
        PORT
        LAYER M3 ;
        RECT  27.840 249.580 28.570 250.000 ;
        LAYER M2 ;
        RECT  27.840 249.580 28.570 250.000 ;
        END
    END I
    PIN VSSO
        DIRECTION INOUT ;
        USE ground ;
        PORT
        LAYER M3 ;
        RECT  0.000 92.060 65.000 123.250 ;
        RECT  64.200 149.940 65.000 162.610 ;
        RECT  0.000 149.940 0.800 162.610 ;
        LAYER M2 ;
        RECT  0.000 147.040 65.000 154.520 ;
        LAYER TOP_M ;
        RECT  0.000 92.060 65.000 123.250 ;
        RECT  0.000 155.410 65.000 162.610 ;
        END
    END VSSO
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        PORT
        LAYER M3 ;
        RECT  64.200 130.690 65.000 148.880 ;
        RECT  0.000 130.690 0.800 148.880 ;
        LAYER M2 ;
        RECT  0.000 136.310 65.000 146.340 ;
        LAYER TOP_M ;
        RECT  0.000 123.850 65.000 154.560 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        PORT
        LAYER M3 ;
        RECT  64.200 163.510 65.000 190.890 ;
        RECT  0.000 163.510 0.800 190.890 ;
        LAYER M2 ;
        RECT  0.000 172.080 65.000 183.060 ;
        LAYER TOP_M ;
        RECT  0.000 163.500 65.000 194.560 ;
        END
    END VDD
    PIN VDDO
        DIRECTION INOUT ;
        USE power ;
        PORT
        LAYER M3 ;
        RECT  64.200 192.330 65.000 200.640 ;
        RECT  0.000 201.660 65.000 221.520 ;
        RECT  0.000 222.720 65.000 246.820 ;
        RECT  0.000 192.330 0.800 200.640 ;
        LAYER M2 ;
        RECT  0.000 186.470 65.000 195.650 ;
        LAYER TOP_M ;
        RECT  0.000 195.170 65.000 200.640 ;
        RECT  0.000 201.660 65.000 221.520 ;
        RECT  0.000 222.720 65.000 246.820 ;
        END
    END VDDO
    OBS
        LAYER M1 ;
        RECT  2.000 0.000 63.000 250.000 ;
        RECT  0.000 88.990 65.000 130.360 ;
        RECT  0.000 136.510 65.000 157.550 ;
        RECT  0.315 158.150 64.700 158.460 ;
        RECT  0.300 158.930 64.700 159.230 ;
        RECT  0.300 159.530 64.700 159.830 ;
        RECT  0.300 160.130 64.700 160.430 ;
        RECT  0.300 160.730 64.700 161.030 ;
        RECT  0.300 161.330 64.700 161.630 ;
        RECT  0.300 161.910 64.700 162.190 ;
        RECT  0.300 162.490 64.700 162.770 ;
        RECT  0.300 163.070 64.700 163.350 ;
        RECT  0.300 163.650 64.700 163.950 ;
        RECT  0.300 164.250 64.700 164.550 ;
        RECT  0.300 164.850 64.700 165.150 ;
        RECT  0.300 165.450 64.700 165.750 ;
        RECT  0.300 166.050 64.700 166.350 ;
        RECT  0.300 166.650 64.700 166.960 ;
        RECT  0.300 167.260 64.700 167.560 ;
        RECT  0.300 167.860 64.700 168.160 ;
        RECT  0.000 169.150 65.000 197.240 ;
        RECT  0.600 0.600 64.400 250.000 ;
        RECT  0.000 198.470 65.000 250.000 ;
        LAYER M2 ;
        RECT  1.840 196.420 2.120 249.400 ;
        RECT  63.180 196.430 63.670 249.400 ;
        RECT  0.600 196.440 64.400 245.485 ;
        RECT  26.530 196.440 64.400 248.790 ;
        RECT  0.600 196.440 22.950 249.400 ;
        RECT  26.530 196.440 27.050 249.400 ;
        RECT  31.420 196.440 64.400 249.400 ;
        RECT  19.140 183.720 52.180 185.680 ;
        RECT  0.600 183.850 64.400 185.680 ;
        RECT  55.195 183.850 56.950 185.850 ;
        RECT  46.230 183.720 51.730 185.870 ;
        RECT  4.830 155.120 7.380 171.290 ;
        RECT  8.170 155.125 8.490 171.290 ;
        RECT  22.160 155.160 22.510 171.290 ;
        RECT  22.810 155.140 23.130 171.290 ;
        RECT  49.290 155.130 51.530 171.290 ;
        RECT  52.470 155.300 52.780 171.290 ;
        RECT  53.655 155.035 53.935 171.290 ;
        RECT  56.365 155.280 56.645 171.315 ;
        RECT  57.120 155.300 57.400 171.315 ;
        RECT  57.835 155.130 58.115 171.315 ;
        RECT  0.600 155.310 64.400 171.290 ;
        RECT  56.240 155.310 61.880 171.315 ;
        RECT  53.895 155.310 55.870 171.370 ;
        RECT  3.175 155.310 3.455 171.380 ;
        RECT  34.655 155.310 38.715 171.480 ;
        RECT  39.605 155.310 42.020 171.480 ;
        RECT  2.000 0.000 63.000 60.210 ;
        RECT  0.600 0.600 64.400 60.210 ;
        RECT  0.600 0.600 1.210 135.520 ;
        RECT  0.600 91.020 64.400 135.520 ;
        RECT  4.080 91.020 60.940 135.690 ;
        RECT  62.580 91.020 62.995 135.710 ;
        LAYER M3 ;
        RECT  0.600 247.660 23.220 248.740 ;
        RECT  0.600 247.660 22.900 249.400 ;
        RECT  26.260 247.660 64.400 248.740 ;
        RECT  26.580 247.660 27.000 249.400 ;
        RECT  31.470 247.660 64.400 249.400 ;
        RECT  0.600 124.090 64.400 129.850 ;
        RECT  1.640 124.090 63.600 135.790 ;
        RECT  1.810 124.090 2.830 154.520 ;
        RECT  3.195 124.090 63.600 171.560 ;
        RECT  3.325 123.900 61.330 171.560 ;
        RECT  1.640 155.040 63.600 171.560 ;
        RECT  1.640 183.580 63.600 185.950 ;
        RECT  5.515 124.090 63.600 200.820 ;
        RECT  1.640 196.170 63.600 200.820 ;
        RECT  56.300 123.900 56.580 201.060 ;
        RECT  0.600 0.600 64.400 60.480 ;
        RECT  2.000 0.000 63.000 88.700 ;
        RECT  0.600 0.600 1.480 91.220 ;
        RECT  0.600 90.750 64.400 91.220 ;
        LAYER TOP_M ;
        RECT  0.600 247.690 64.400 248.850 ;
        RECT  0.600 247.690 23.010 249.400 ;
        RECT  26.470 247.690 27.110 249.400 ;
        RECT  31.360 247.690 64.400 249.400 ;
        RECT  2.000 0.000 63.000 91.190 ;
        RECT  0.600 0.600 64.400 91.190 ;
    END
END pc3b04d

MACRO pc3b04
    CLASS PAD ;
    FOREIGN pc3b04 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 65.000 BY 250.000 ;
    SYMMETRY X Y R90 ;
    SITE IOSite_c ;
    PIN PAD
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 55.440  LAYER TOP_M  ;
        ANTENNAPARTIALMETALSIDEAREA 287.938  LAYER M3  ;
        ANTENNAPARTIALMETALSIDEAREA 480.740  LAYER M2  ;
        ANTENNADIFFAREA 2657.280  LAYER TOP_M  ;
        ANTENNADIFFAREA 1209.600  LAYER M2  ;
        ANTENNADIFFAREA 2657.280  LAYER M3  ;
        ANTENNAPARTIALCUTAREA 632.318  LAYER TOP_V  ;
        ANTENNAPARTIALCUTAREA 349.898  LAYER V3  ;
        ANTENNAPARTIALCUTAREA 255.798  LAYER V2  ;
        PORT
        LAYER M3 ;
        RECT  23.740 249.580 25.740 250.000 ;
        LAYER M2 ;
        RECT  2.000 61.000 63.000 90.230 ;
        RECT  23.740 246.275 25.740 250.000 ;
        END
    END PAD
    PIN OEN
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 80.634  LAYER M2  ;
        ANTENNAPARTIALMETALSIDEAREA 41.679  LAYER M3  ;
        ANTENNAPARTIALMETALSIDEAREA 67.374  LAYER M1  ;
        ANTENNADIFFAREA 0.250  LAYER M3  ;
        ANTENNAPARTIALCUTAREA 0.203  LAYER V2  ;
        ANTENNAPARTIALCUTAREA 0.135  LAYER V3  ;
        ANTENNAGATEAREA 9.900  LAYER M3  ;
        ANTENNAGATEAREA 8.100  LAYER M2  ;
        PORT
        LAYER M3 ;
        RECT  29.900 249.580 30.630 250.000 ;
        LAYER M2 ;
        RECT  29.900 249.580 30.630 250.000 ;
        END
    END OEN
    PIN CIN
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 32.277  LAYER M3  ;
        ANTENNAPARTIALMETALSIDEAREA 96.916  LAYER M2  ;
        ANTENNAPARTIALMETALSIDEAREA 67.374  LAYER M1  ;
        ANTENNADIFFAREA 20.600  LAYER M3  ;
        ANTENNAPARTIALCUTAREA 0.135  LAYER V3  ;
        ANTENNAPARTIALCUTAREA 0.203  LAYER V2  ;
        PORT
        LAYER M3 ;
        RECT  28.870 249.580 29.600 250.000 ;
        LAYER M2 ;
        RECT  28.870 249.580 29.600 250.000 ;
        END
    END CIN
    PIN I
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 67.374  LAYER M1  ;
        ANTENNAPARTIALMETALSIDEAREA 80.804  LAYER M2  ;
        ANTENNAPARTIALMETALSIDEAREA 41.096  LAYER M3  ;
        ANTENNADIFFAREA 0.250  LAYER M3  ;
        ANTENNAPARTIALCUTAREA 0.270  LAYER V2  ;
        ANTENNAPARTIALCUTAREA 0.135  LAYER V3  ;
        ANTENNAGATEAREA 18.900  LAYER M2  ;
        ANTENNAGATEAREA 20.700  LAYER M3  ;
        PORT
        LAYER M3 ;
        RECT  27.840 249.580 28.570 250.000 ;
        LAYER M2 ;
        RECT  27.840 249.580 28.570 250.000 ;
        END
    END I
    PIN VSSO
        DIRECTION INOUT ;
        USE ground ;
        PORT
        LAYER M3 ;
        RECT  0.000 92.060 65.000 123.250 ;
        RECT  64.200 149.940 65.000 162.610 ;
        RECT  0.000 149.940 0.800 162.610 ;
        LAYER M2 ;
        RECT  0.000 147.040 65.000 154.520 ;
        LAYER TOP_M ;
        RECT  0.000 92.060 65.000 123.250 ;
        RECT  0.000 155.410 65.000 162.610 ;
        END
    END VSSO
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        PORT
        LAYER M3 ;
        RECT  64.200 130.690 65.000 148.880 ;
        RECT  0.000 130.690 0.800 148.880 ;
        LAYER M2 ;
        RECT  0.000 136.310 65.000 146.340 ;
        LAYER TOP_M ;
        RECT  0.000 123.850 65.000 154.560 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        PORT
        LAYER M3 ;
        RECT  64.200 163.510 65.000 190.890 ;
        RECT  0.000 163.510 0.800 190.890 ;
        LAYER M2 ;
        RECT  0.000 172.080 65.000 183.060 ;
        LAYER TOP_M ;
        RECT  0.000 163.500 65.000 194.560 ;
        END
    END VDD
    PIN VDDO
        DIRECTION INOUT ;
        USE power ;
        PORT
        LAYER M3 ;
        RECT  64.200 192.330 65.000 200.640 ;
        RECT  0.000 201.660 65.000 221.520 ;
        RECT  0.000 222.720 65.000 246.820 ;
        RECT  0.000 192.330 0.800 200.640 ;
        LAYER M2 ;
        RECT  0.000 186.470 65.000 195.650 ;
        LAYER TOP_M ;
        RECT  0.000 195.170 65.000 200.640 ;
        RECT  0.000 201.660 65.000 221.520 ;
        RECT  0.000 222.720 65.000 246.820 ;
        END
    END VDDO
    OBS
        LAYER M1 ;
        RECT  2.000 0.000 63.000 250.000 ;
        RECT  0.000 88.990 65.000 130.360 ;
        RECT  0.000 136.510 65.000 157.550 ;
        RECT  0.315 158.150 64.700 158.460 ;
        RECT  0.300 158.930 64.700 159.230 ;
        RECT  0.300 159.530 64.700 159.830 ;
        RECT  0.300 160.130 64.700 160.430 ;
        RECT  0.300 160.730 64.700 161.030 ;
        RECT  0.300 161.330 64.700 161.630 ;
        RECT  0.300 161.910 64.700 162.190 ;
        RECT  0.300 162.490 64.700 162.770 ;
        RECT  0.300 163.070 64.700 163.350 ;
        RECT  0.300 163.650 64.700 163.950 ;
        RECT  0.300 164.250 64.700 164.550 ;
        RECT  0.300 164.850 64.700 165.150 ;
        RECT  0.300 165.450 64.700 165.750 ;
        RECT  0.300 166.050 64.700 166.350 ;
        RECT  0.300 166.650 64.700 166.960 ;
        RECT  0.300 167.260 64.700 167.560 ;
        RECT  0.300 167.860 64.700 168.160 ;
        RECT  0.000 169.150 65.000 197.240 ;
        RECT  0.600 0.600 64.400 250.000 ;
        RECT  0.000 198.470 65.000 250.000 ;
        LAYER M2 ;
        RECT  1.840 196.420 2.120 249.400 ;
        RECT  63.180 196.430 63.670 249.400 ;
        RECT  0.600 196.440 64.400 245.485 ;
        RECT  26.530 196.440 64.400 248.790 ;
        RECT  0.600 196.440 22.950 249.400 ;
        RECT  26.530 196.440 27.050 249.400 ;
        RECT  31.420 196.440 64.400 249.400 ;
        RECT  19.140 183.720 52.180 185.680 ;
        RECT  0.600 183.850 64.400 185.680 ;
        RECT  55.195 183.850 56.950 185.850 ;
        RECT  46.230 183.720 51.730 185.870 ;
        RECT  4.830 155.120 7.380 171.290 ;
        RECT  8.170 155.125 8.490 171.290 ;
        RECT  22.160 155.160 22.510 171.290 ;
        RECT  22.810 155.140 23.130 171.290 ;
        RECT  53.655 155.035 53.935 171.290 ;
        RECT  56.365 155.280 56.645 171.315 ;
        RECT  57.120 155.300 57.400 171.315 ;
        RECT  57.835 155.130 58.115 171.315 ;
        RECT  0.600 155.310 64.400 171.290 ;
        RECT  56.240 155.310 61.880 171.315 ;
        RECT  53.895 155.310 55.870 171.370 ;
        RECT  3.175 155.310 3.455 171.380 ;
        RECT  34.655 155.310 38.715 171.480 ;
        RECT  39.605 155.310 42.020 171.480 ;
        RECT  2.000 0.000 63.000 60.210 ;
        RECT  0.600 0.600 64.400 60.210 ;
        RECT  0.600 0.600 1.210 135.520 ;
        RECT  0.600 91.020 64.400 135.520 ;
        RECT  4.080 91.020 60.940 135.690 ;
        RECT  62.580 91.020 62.995 135.710 ;
        LAYER M3 ;
        RECT  0.600 247.660 23.220 248.740 ;
        RECT  0.600 247.660 22.900 249.400 ;
        RECT  26.260 247.660 64.400 248.740 ;
        RECT  26.580 247.660 27.000 249.400 ;
        RECT  31.470 247.660 64.400 249.400 ;
        RECT  0.600 124.090 64.400 129.850 ;
        RECT  1.640 124.090 63.600 135.790 ;
        RECT  1.810 124.090 2.830 154.520 ;
        RECT  3.195 124.090 63.600 171.560 ;
        RECT  3.325 123.900 61.330 171.560 ;
        RECT  1.640 155.040 63.600 171.560 ;
        RECT  1.640 183.580 63.600 185.950 ;
        RECT  5.515 124.090 63.600 200.820 ;
        RECT  1.640 196.170 63.600 200.820 ;
        RECT  56.300 123.900 56.580 201.060 ;
        RECT  0.600 0.600 64.400 60.480 ;
        RECT  2.000 0.000 63.000 88.700 ;
        RECT  0.600 0.600 1.480 91.220 ;
        RECT  0.600 90.750 64.400 91.220 ;
        LAYER TOP_M ;
        RECT  0.600 247.690 64.400 248.850 ;
        RECT  0.600 247.690 23.010 249.400 ;
        RECT  26.470 247.690 27.110 249.400 ;
        RECT  31.360 247.690 64.400 249.400 ;
        RECT  2.000 0.000 63.000 91.190 ;
        RECT  0.600 0.600 64.400 91.190 ;
    END
END pc3b04

MACRO pc3b03u
    CLASS PAD ;
    FOREIGN pc3b03u 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 65.000 BY 250.000 ;
    SYMMETRY X Y R90 ;
    SITE IOSite_c ;
    PIN PAD
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 55.440  LAYER TOP_M  ;
        ANTENNAPARTIALMETALSIDEAREA 287.938  LAYER M3  ;
        ANTENNAPARTIALMETALSIDEAREA 480.740  LAYER M2  ;
        ANTENNADIFFAREA 2657.280  LAYER TOP_M  ;
        ANTENNADIFFAREA 1209.600  LAYER M2  ;
        ANTENNADIFFAREA 2657.280  LAYER M3  ;
        ANTENNAPARTIALCUTAREA 632.318  LAYER TOP_V  ;
        ANTENNAPARTIALCUTAREA 349.898  LAYER V3  ;
        ANTENNAPARTIALCUTAREA 255.798  LAYER V2  ;
        PORT
        LAYER M3 ;
        RECT  23.740 249.580 25.740 250.000 ;
        LAYER M2 ;
        RECT  2.000 61.000 63.000 90.230 ;
        RECT  23.740 246.275 25.740 250.000 ;
        END
    END PAD
    PIN OEN
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 80.634  LAYER M2  ;
        ANTENNAPARTIALMETALSIDEAREA 41.679  LAYER M3  ;
        ANTENNAPARTIALMETALSIDEAREA 67.374  LAYER M1  ;
        ANTENNADIFFAREA 0.250  LAYER M3  ;
        ANTENNAPARTIALCUTAREA 0.203  LAYER V2  ;
        ANTENNAPARTIALCUTAREA 0.135  LAYER V3  ;
        ANTENNAGATEAREA 9.900  LAYER M3  ;
        ANTENNAGATEAREA 8.100  LAYER M2  ;
        PORT
        LAYER M3 ;
        RECT  29.900 249.580 30.630 250.000 ;
        LAYER M2 ;
        RECT  29.900 249.580 30.630 250.000 ;
        END
    END OEN
    PIN CIN
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 32.277  LAYER M3  ;
        ANTENNAPARTIALMETALSIDEAREA 96.916  LAYER M2  ;
        ANTENNAPARTIALMETALSIDEAREA 67.374  LAYER M1  ;
        ANTENNADIFFAREA 20.600  LAYER M3  ;
        ANTENNAPARTIALCUTAREA 0.135  LAYER V3  ;
        ANTENNAPARTIALCUTAREA 0.203  LAYER V2  ;
        PORT
        LAYER M3 ;
        RECT  28.870 249.580 29.600 250.000 ;
        LAYER M2 ;
        RECT  28.870 249.580 29.600 250.000 ;
        END
    END CIN
    PIN I
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 67.374  LAYER M1  ;
        ANTENNAPARTIALMETALSIDEAREA 80.804  LAYER M2  ;
        ANTENNAPARTIALMETALSIDEAREA 41.096  LAYER M3  ;
        ANTENNADIFFAREA 0.250  LAYER M3  ;
        ANTENNAPARTIALCUTAREA 0.270  LAYER V2  ;
        ANTENNAPARTIALCUTAREA 0.135  LAYER V3  ;
        ANTENNAGATEAREA 18.900  LAYER M2  ;
        ANTENNAGATEAREA 20.700  LAYER M3  ;
        PORT
        LAYER M3 ;
        RECT  27.840 249.580 28.570 250.000 ;
        LAYER M2 ;
        RECT  27.840 249.580 28.570 250.000 ;
        END
    END I
    PIN VDDO
        DIRECTION INOUT ;
        USE power ;
        PORT
        LAYER M3 ;
        RECT  64.200 192.330 65.000 200.640 ;
        RECT  0.000 201.660 65.000 221.520 ;
        RECT  0.000 222.720 65.000 246.820 ;
        RECT  0.000 192.330 0.800 200.640 ;
        LAYER M2 ;
        RECT  0.000 186.470 65.000 195.650 ;
        LAYER TOP_M ;
        RECT  0.000 195.170 65.000 200.640 ;
        RECT  0.000 201.660 65.000 221.520 ;
        RECT  0.000 222.720 65.000 246.820 ;
        END
    END VDDO
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        PORT
        LAYER M3 ;
        RECT  64.200 163.510 65.000 190.890 ;
        RECT  0.000 163.510 0.800 190.890 ;
        LAYER M2 ;
        RECT  0.000 172.080 65.000 183.060 ;
        LAYER TOP_M ;
        RECT  0.000 163.500 65.000 194.560 ;
        END
    END VDD
    PIN VSSO
        DIRECTION INOUT ;
        USE ground ;
        PORT
        LAYER M3 ;
        RECT  0.000 92.060 65.000 123.250 ;
        RECT  64.200 149.940 65.000 162.610 ;
        RECT  0.000 149.940 0.800 162.610 ;
        LAYER M2 ;
        RECT  0.000 147.040 65.000 154.520 ;
        LAYER TOP_M ;
        RECT  0.000 92.060 65.000 123.250 ;
        RECT  0.000 155.410 65.000 162.610 ;
        END
    END VSSO
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        PORT
        LAYER M3 ;
        RECT  64.200 130.690 65.000 148.880 ;
        RECT  0.000 130.690 0.800 148.880 ;
        LAYER M2 ;
        RECT  0.000 136.310 65.000 146.340 ;
        LAYER TOP_M ;
        RECT  0.000 123.850 65.000 154.560 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  2.000 0.000 63.000 250.000 ;
        RECT  0.000 88.990 65.000 130.360 ;
        RECT  0.000 136.510 65.000 157.550 ;
        RECT  0.315 158.150 64.700 158.460 ;
        RECT  0.300 158.930 64.700 159.230 ;
        RECT  0.300 159.530 64.700 159.830 ;
        RECT  0.300 160.130 64.700 160.430 ;
        RECT  0.300 160.730 64.700 161.030 ;
        RECT  0.300 161.330 64.700 161.630 ;
        RECT  0.300 161.910 64.700 162.190 ;
        RECT  0.300 162.490 64.700 162.770 ;
        RECT  0.300 163.070 64.700 163.350 ;
        RECT  0.300 163.650 64.700 163.950 ;
        RECT  0.300 164.250 64.700 164.550 ;
        RECT  0.300 164.850 64.700 165.150 ;
        RECT  0.300 165.450 64.700 165.750 ;
        RECT  0.300 166.050 64.700 166.350 ;
        RECT  0.300 166.650 64.700 166.960 ;
        RECT  0.300 167.260 64.700 167.560 ;
        RECT  0.300 167.860 64.700 168.160 ;
        RECT  0.000 169.150 65.000 197.240 ;
        RECT  0.600 0.600 64.400 250.000 ;
        RECT  0.000 198.470 65.000 250.000 ;
        LAYER M2 ;
        RECT  1.840 196.420 2.120 249.400 ;
        RECT  63.180 196.430 63.670 249.400 ;
        RECT  0.600 196.440 64.400 245.485 ;
        RECT  26.530 196.440 64.400 248.790 ;
        RECT  0.600 196.440 22.950 249.400 ;
        RECT  26.530 196.440 27.050 249.400 ;
        RECT  31.420 196.440 64.400 249.400 ;
        RECT  19.440 183.720 52.185 185.680 ;
        RECT  0.600 183.850 64.400 185.680 ;
        RECT  46.230 183.720 51.730 185.870 ;
        RECT  54.855 183.850 56.700 185.950 ;
        RECT  4.895 155.120 7.525 171.290 ;
        RECT  8.170 155.125 8.490 171.290 ;
        RECT  22.160 155.160 22.510 171.290 ;
        RECT  22.810 155.140 23.130 171.290 ;
        RECT  53.655 155.035 53.935 171.290 ;
        RECT  56.365 155.280 56.645 171.315 ;
        RECT  57.120 155.300 57.400 171.315 ;
        RECT  57.835 155.130 58.115 171.315 ;
        RECT  0.600 155.310 64.400 171.290 ;
        RECT  56.240 155.310 61.880 171.315 ;
        RECT  33.625 155.310 34.125 171.365 ;
        RECT  53.895 155.310 55.870 171.370 ;
        RECT  3.220 155.310 3.500 171.380 ;
        RECT  34.655 155.310 38.715 171.480 ;
        RECT  39.605 155.310 42.020 171.480 ;
        RECT  2.000 0.000 63.000 60.210 ;
        RECT  0.600 0.600 64.400 60.210 ;
        RECT  0.600 0.600 1.210 135.520 ;
        RECT  0.600 91.020 64.400 135.520 ;
        RECT  4.080 91.020 60.940 135.690 ;
        RECT  62.580 91.020 62.995 135.710 ;
        LAYER M3 ;
        RECT  0.600 247.660 23.220 248.740 ;
        RECT  0.600 247.660 22.900 249.400 ;
        RECT  26.260 247.660 64.400 248.740 ;
        RECT  26.580 247.660 27.000 249.400 ;
        RECT  31.470 247.660 64.400 249.400 ;
        RECT  0.600 124.090 64.400 129.850 ;
        RECT  1.640 124.090 63.600 135.790 ;
        RECT  1.810 124.090 2.830 154.520 ;
        RECT  3.110 124.090 63.600 171.560 ;
        RECT  4.040 123.970 60.900 171.560 ;
        RECT  1.640 155.040 63.600 171.560 ;
        RECT  1.640 183.580 63.600 185.950 ;
        RECT  5.510 124.090 63.600 200.820 ;
        RECT  1.640 196.170 63.600 200.820 ;
        RECT  56.300 123.970 56.580 201.060 ;
        RECT  0.600 0.600 64.400 60.480 ;
        RECT  2.000 0.000 63.000 88.700 ;
        RECT  0.600 0.600 1.480 91.220 ;
        RECT  0.600 90.750 64.400 91.220 ;
        LAYER TOP_M ;
        RECT  0.600 247.690 64.400 248.850 ;
        RECT  0.600 247.690 23.010 249.400 ;
        RECT  26.470 247.690 27.110 249.400 ;
        RECT  31.360 247.690 64.400 249.400 ;
        RECT  2.000 0.000 63.000 91.190 ;
        RECT  0.600 0.600 64.400 91.190 ;
    END
END pc3b03u

MACRO pc3b03ed
    CLASS PAD ;
    FOREIGN pc3b03ed 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 65.000 BY 250.000 ;
    SYMMETRY X Y R90 ;
    SITE IOSite_c ;
    PIN RENB
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 82.012  LAYER M2  ;
        ANTENNAPARTIALMETALSIDEAREA 44.266  LAYER M3  ;
        ANTENNADIFFAREA 1.000  LAYER M3  ;
        ANTENNAPARTIALCUTAREA 0.135  LAYER V3  ;
        ANTENNAGATEAREA 6.316  LAYER M3  ;
        PORT
        LAYER M3 ;
        RECT  30.930 249.580 31.660 250.000 ;
        LAYER M2 ;
        RECT  30.930 249.580 31.660 250.000 ;
        END
    END RENB
    PIN PAD
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 55.440  LAYER TOP_M  ;
        ANTENNAPARTIALMETALSIDEAREA 287.938  LAYER M3  ;
        ANTENNAPARTIALMETALSIDEAREA 480.740  LAYER M2  ;
        ANTENNADIFFAREA 2657.280  LAYER TOP_M  ;
        ANTENNADIFFAREA 2657.280  LAYER M3  ;
        ANTENNADIFFAREA 1209.600  LAYER M2  ;
        ANTENNAPARTIALCUTAREA 632.318  LAYER TOP_V  ;
        ANTENNAPARTIALCUTAREA 349.898  LAYER V3  ;
        ANTENNAPARTIALCUTAREA 255.798  LAYER V2  ;
        PORT
        LAYER M3 ;
        RECT  23.740 249.580 25.740 250.000 ;
        LAYER M2 ;
        RECT  2.000 61.000 63.000 90.230 ;
        RECT  23.740 246.275 25.740 250.000 ;
        END
    END PAD
    PIN OEN
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 67.480  LAYER M3  ;
        ANTENNAPARTIALMETALSIDEAREA 79.336  LAYER M2  ;
        ANTENNAPARTIALMETALSIDEAREA 67.374  LAYER M1  ;
        ANTENNADIFFAREA 0.250  LAYER M3  ;
        ANTENNAPARTIALCUTAREA 0.135  LAYER V3  ;
        ANTENNAPARTIALCUTAREA 0.338  LAYER V2  ;
        ANTENNAGATEAREA 8.100  LAYER M2  ;
        ANTENNAGATEAREA 9.900  LAYER M3  ;
        PORT
        LAYER M3 ;
        RECT  29.900 249.580 30.630 250.000 ;
        LAYER M2 ;
        RECT  29.900 249.580 30.630 250.000 ;
        END
    END OEN
    PIN CIN
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 67.374  LAYER M1  ;
        ANTENNAPARTIALMETALSIDEAREA 79.134  LAYER M2  ;
        ANTENNAPARTIALMETALSIDEAREA 40.964  LAYER M3  ;
        ANTENNADIFFAREA 20.727  LAYER M3  ;
        ANTENNAPARTIALCUTAREA 0.135  LAYER V3  ;
        ANTENNAPARTIALCUTAREA 0.203  LAYER V2  ;
        PORT
        LAYER M3 ;
        RECT  28.870 249.580 29.600 250.000 ;
        LAYER M2 ;
        RECT  28.870 249.580 29.600 250.000 ;
        END
    END CIN
    PIN I
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 67.374  LAYER M1  ;
        ANTENNAPARTIALMETALSIDEAREA 79.415  LAYER M2  ;
        ANTENNAPARTIALMETALSIDEAREA 42.050  LAYER M3  ;
        ANTENNADIFFAREA 0.250  LAYER M3  ;
        ANTENNAPARTIALCUTAREA 0.270  LAYER V2  ;
        ANTENNAPARTIALCUTAREA 0.135  LAYER V3  ;
        ANTENNAGATEAREA 18.900  LAYER M2  ;
        ANTENNAGATEAREA 20.700  LAYER M3  ;
        PORT
        LAYER M3 ;
        RECT  27.840 249.580 28.570 250.000 ;
        LAYER M2 ;
        RECT  27.840 249.580 28.570 250.000 ;
        END
    END I
    PIN VDDO
        DIRECTION INOUT ;
        USE power ;
        PORT
        LAYER M3 ;
        RECT  64.200 192.330 65.000 200.640 ;
        RECT  0.000 201.660 65.000 221.520 ;
        RECT  0.000 222.720 65.000 246.820 ;
        RECT  0.000 192.330 0.800 200.640 ;
        LAYER M2 ;
        RECT  0.000 186.470 65.000 195.650 ;
        LAYER TOP_M ;
        RECT  0.000 195.170 65.000 200.640 ;
        RECT  0.000 201.660 65.000 221.520 ;
        RECT  0.000 222.720 65.000 246.820 ;
        END
    END VDDO
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        PORT
        LAYER M3 ;
        RECT  64.200 163.510 65.000 190.890 ;
        RECT  0.000 163.510 0.800 190.890 ;
        LAYER M2 ;
        RECT  0.000 172.080 65.000 183.060 ;
        LAYER TOP_M ;
        RECT  0.000 163.500 65.000 194.560 ;
        END
    END VDD
    PIN VSSO
        DIRECTION INOUT ;
        USE ground ;
        PORT
        LAYER M3 ;
        RECT  0.000 92.060 65.000 123.250 ;
        RECT  64.200 149.940 65.000 162.610 ;
        RECT  0.000 149.940 0.800 162.610 ;
        LAYER M2 ;
        RECT  0.000 147.040 65.000 154.520 ;
        LAYER TOP_M ;
        RECT  0.000 92.060 65.000 123.250 ;
        RECT  0.000 155.410 65.000 162.610 ;
        END
    END VSSO
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        PORT
        LAYER M3 ;
        RECT  64.200 130.690 65.000 148.880 ;
        RECT  0.000 130.690 0.800 148.880 ;
        LAYER M2 ;
        RECT  0.000 136.310 65.000 146.340 ;
        LAYER TOP_M ;
        RECT  0.000 123.850 65.000 154.560 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  2.000 0.000 63.000 250.000 ;
        RECT  0.000 88.990 65.000 130.360 ;
        RECT  0.000 136.510 65.000 157.550 ;
        RECT  0.300 158.330 64.700 158.630 ;
        RECT  0.300 158.930 64.700 159.230 ;
        RECT  0.300 159.530 64.700 159.830 ;
        RECT  0.300 160.130 64.700 160.430 ;
        RECT  0.300 160.730 64.700 161.030 ;
        RECT  0.300 161.330 64.700 161.630 ;
        RECT  0.300 161.910 64.700 162.190 ;
        RECT  0.300 162.490 64.700 162.770 ;
        RECT  0.300 163.070 64.700 163.350 ;
        RECT  0.300 163.650 64.700 163.950 ;
        RECT  0.300 164.250 64.700 164.550 ;
        RECT  0.300 164.850 64.700 165.150 ;
        RECT  0.300 165.450 64.700 165.750 ;
        RECT  0.300 166.050 64.700 166.350 ;
        RECT  0.300 166.650 64.700 166.960 ;
        RECT  0.300 167.260 64.700 167.560 ;
        RECT  0.300 167.860 64.700 168.160 ;
        RECT  0.000 169.150 65.000 197.240 ;
        RECT  0.600 0.600 64.400 250.000 ;
        RECT  0.000 198.470 65.000 250.000 ;
        LAYER M2 ;
        RECT  1.740 196.420 2.020 249.400 ;
        RECT  63.180 196.430 63.670 249.400 ;
        RECT  0.600 196.440 64.400 245.485 ;
        RECT  26.530 196.440 64.400 248.790 ;
        RECT  0.600 196.440 22.950 249.400 ;
        RECT  26.530 196.440 27.050 249.400 ;
        RECT  32.450 196.440 64.400 249.400 ;
        RECT  19.440 183.720 52.185 185.680 ;
        RECT  55.995 183.710 56.315 185.880 ;
        RECT  0.600 183.850 64.400 185.680 ;
        RECT  46.230 183.720 51.730 185.870 ;
        RECT  54.085 183.850 54.915 185.870 ;
        RECT  55.375 183.850 61.350 185.880 ;
        RECT  4.895 155.120 7.525 171.290 ;
        RECT  8.170 155.125 8.490 171.290 ;
        RECT  22.160 155.160 22.510 171.290 ;
        RECT  22.810 155.140 23.130 171.290 ;
        RECT  32.135 155.120 32.415 171.290 ;
        RECT  32.695 155.120 34.425 171.290 ;
        RECT  48.835 155.120 49.155 171.290 ;
        RECT  49.535 155.120 49.815 171.290 ;
        RECT  50.120 155.125 50.450 171.290 ;
        RECT  51.785 155.120 53.330 171.290 ;
        RECT  53.695 155.110 53.995 171.325 ;
        RECT  57.755 155.130 58.035 171.290 ;
        RECT  0.600 155.310 64.400 171.290 ;
        RECT  15.415 155.310 15.915 171.295 ;
        RECT  53.055 155.310 57.850 171.325 ;
        RECT  3.220 155.310 3.500 171.380 ;
        RECT  33.355 155.310 39.260 171.480 ;
        RECT  41.105 155.310 43.490 171.480 ;
        RECT  60.240 155.310 63.080 171.480 ;
        RECT  2.000 0.000 63.000 60.210 ;
        RECT  0.600 0.600 64.400 60.210 ;
        RECT  0.600 0.600 1.210 135.520 ;
        RECT  0.600 91.020 64.400 135.520 ;
        RECT  4.080 91.020 60.940 135.690 ;
        RECT  62.580 91.020 62.995 135.710 ;
        LAYER M3 ;
        RECT  0.600 247.660 23.220 248.740 ;
        RECT  0.600 247.660 22.900 249.400 ;
        RECT  26.260 247.660 64.400 248.740 ;
        RECT  26.580 247.660 27.000 249.400 ;
        RECT  32.500 247.660 64.400 249.400 ;
        RECT  0.600 124.090 64.400 129.850 ;
        RECT  1.640 124.090 63.600 135.790 ;
        RECT  1.810 124.090 2.830 154.520 ;
        RECT  3.110 124.090 63.600 171.560 ;
        RECT  4.040 123.970 60.900 171.560 ;
        RECT  1.640 155.040 63.600 171.560 ;
        RECT  1.640 183.580 63.600 185.950 ;
        RECT  5.510 124.090 63.600 200.820 ;
        RECT  1.640 196.170 63.600 200.820 ;
        RECT  54.265 123.970 54.545 201.060 ;
        RECT  0.600 0.600 64.400 60.480 ;
        RECT  2.000 0.000 63.000 88.700 ;
        RECT  0.600 0.600 1.480 91.220 ;
        RECT  0.600 90.750 64.400 91.220 ;
        LAYER TOP_M ;
        RECT  0.600 247.690 64.400 248.850 ;
        RECT  0.600 247.690 23.010 249.400 ;
        RECT  26.470 247.690 27.110 249.400 ;
        RECT  32.390 247.690 64.400 249.400 ;
        RECT  2.000 0.000 63.000 91.190 ;
        RECT  0.600 0.600 64.400 91.190 ;
    END
END pc3b03ed

MACRO pc3b03d
    CLASS PAD ;
    FOREIGN pc3b03d 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 65.000 BY 250.000 ;
    SYMMETRY X Y R90 ;
    SITE IOSite_c ;
    PIN PAD
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 55.440  LAYER TOP_M  ;
        ANTENNAPARTIALMETALSIDEAREA 287.938  LAYER M3  ;
        ANTENNAPARTIALMETALSIDEAREA 480.740  LAYER M2  ;
        ANTENNADIFFAREA 2657.280  LAYER TOP_M  ;
        ANTENNADIFFAREA 1209.600  LAYER M2  ;
        ANTENNADIFFAREA 2657.280  LAYER M3  ;
        ANTENNAPARTIALCUTAREA 632.318  LAYER TOP_V  ;
        ANTENNAPARTIALCUTAREA 349.898  LAYER V3  ;
        ANTENNAPARTIALCUTAREA 255.798  LAYER V2  ;
        PORT
        LAYER M3 ;
        RECT  23.740 249.580 25.740 250.000 ;
        LAYER M2 ;
        RECT  2.000 61.000 63.000 90.230 ;
        RECT  23.740 246.275 25.740 250.000 ;
        END
    END PAD
    PIN OEN
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 80.634  LAYER M2  ;
        ANTENNAPARTIALMETALSIDEAREA 41.679  LAYER M3  ;
        ANTENNAPARTIALMETALSIDEAREA 67.374  LAYER M1  ;
        ANTENNADIFFAREA 0.250  LAYER M3  ;
        ANTENNAPARTIALCUTAREA 0.203  LAYER V2  ;
        ANTENNAPARTIALCUTAREA 0.135  LAYER V3  ;
        ANTENNAGATEAREA 9.900  LAYER M3  ;
        ANTENNAGATEAREA 8.100  LAYER M2  ;
        PORT
        LAYER M3 ;
        RECT  29.900 249.580 30.630 250.000 ;
        LAYER M2 ;
        RECT  29.900 249.580 30.630 250.000 ;
        END
    END OEN
    PIN CIN
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 32.277  LAYER M3  ;
        ANTENNAPARTIALMETALSIDEAREA 96.916  LAYER M2  ;
        ANTENNAPARTIALMETALSIDEAREA 67.374  LAYER M1  ;
        ANTENNADIFFAREA 20.600  LAYER M3  ;
        ANTENNAPARTIALCUTAREA 0.135  LAYER V3  ;
        ANTENNAPARTIALCUTAREA 0.203  LAYER V2  ;
        PORT
        LAYER M3 ;
        RECT  28.870 249.580 29.600 250.000 ;
        LAYER M2 ;
        RECT  28.870 249.580 29.600 250.000 ;
        END
    END CIN
    PIN I
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 67.374  LAYER M1  ;
        ANTENNAPARTIALMETALSIDEAREA 80.804  LAYER M2  ;
        ANTENNAPARTIALMETALSIDEAREA 41.096  LAYER M3  ;
        ANTENNADIFFAREA 0.250  LAYER M3  ;
        ANTENNAPARTIALCUTAREA 0.270  LAYER V2  ;
        ANTENNAPARTIALCUTAREA 0.135  LAYER V3  ;
        ANTENNAGATEAREA 18.900  LAYER M2  ;
        ANTENNAGATEAREA 20.700  LAYER M3  ;
        PORT
        LAYER M3 ;
        RECT  27.840 249.580 28.570 250.000 ;
        LAYER M2 ;
        RECT  27.840 249.580 28.570 250.000 ;
        END
    END I
    PIN VDDO
        DIRECTION INOUT ;
        USE power ;
        PORT
        LAYER M3 ;
        RECT  64.200 192.330 65.000 200.640 ;
        RECT  0.000 201.660 65.000 221.520 ;
        RECT  0.000 222.720 65.000 246.820 ;
        RECT  0.000 192.330 0.800 200.640 ;
        LAYER M2 ;
        RECT  0.000 186.470 65.000 195.650 ;
        LAYER TOP_M ;
        RECT  0.000 195.170 65.000 200.640 ;
        RECT  0.000 201.660 65.000 221.520 ;
        RECT  0.000 222.720 65.000 246.820 ;
        END
    END VDDO
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        PORT
        LAYER M3 ;
        RECT  64.200 163.510 65.000 190.890 ;
        RECT  0.000 163.510 0.800 190.890 ;
        LAYER M2 ;
        RECT  0.000 172.080 65.000 183.060 ;
        LAYER TOP_M ;
        RECT  0.000 163.500 65.000 194.560 ;
        END
    END VDD
    PIN VSSO
        DIRECTION INOUT ;
        USE ground ;
        PORT
        LAYER M3 ;
        RECT  0.000 92.060 65.000 123.250 ;
        RECT  64.200 149.940 65.000 162.610 ;
        RECT  0.000 149.940 0.800 162.610 ;
        LAYER M2 ;
        RECT  0.000 147.040 65.000 154.520 ;
        LAYER TOP_M ;
        RECT  0.000 92.060 65.000 123.250 ;
        RECT  0.000 155.410 65.000 162.610 ;
        END
    END VSSO
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        PORT
        LAYER M3 ;
        RECT  64.200 130.690 65.000 148.880 ;
        RECT  0.000 130.690 0.800 148.880 ;
        LAYER M2 ;
        RECT  0.000 136.310 65.000 146.340 ;
        LAYER TOP_M ;
        RECT  0.000 123.850 65.000 154.560 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  2.000 0.000 63.000 250.000 ;
        RECT  0.000 88.990 65.000 130.360 ;
        RECT  0.000 136.510 65.000 157.550 ;
        RECT  0.315 158.150 64.700 158.460 ;
        RECT  0.300 158.930 64.700 159.230 ;
        RECT  0.300 159.530 64.700 159.830 ;
        RECT  0.300 160.130 64.700 160.430 ;
        RECT  0.300 160.730 64.700 161.030 ;
        RECT  0.300 161.330 64.700 161.630 ;
        RECT  0.300 161.910 64.700 162.190 ;
        RECT  0.300 162.490 64.700 162.770 ;
        RECT  0.300 163.070 64.700 163.350 ;
        RECT  0.300 163.650 64.700 163.950 ;
        RECT  0.300 164.250 64.700 164.550 ;
        RECT  0.300 164.850 64.700 165.150 ;
        RECT  0.300 165.450 64.700 165.750 ;
        RECT  0.300 166.050 64.700 166.350 ;
        RECT  0.300 166.650 64.700 166.960 ;
        RECT  0.300 167.260 64.700 167.560 ;
        RECT  0.300 167.860 64.700 168.160 ;
        RECT  0.000 169.150 65.000 197.240 ;
        RECT  0.600 0.600 64.400 250.000 ;
        RECT  0.000 198.470 65.000 250.000 ;
        LAYER M2 ;
        RECT  1.840 196.420 2.120 249.400 ;
        RECT  63.180 196.430 63.670 249.400 ;
        RECT  0.600 196.440 64.400 245.485 ;
        RECT  26.530 196.440 64.400 248.790 ;
        RECT  0.600 196.440 22.950 249.400 ;
        RECT  26.530 196.440 27.050 249.400 ;
        RECT  31.420 196.440 64.400 249.400 ;
        RECT  19.440 183.720 52.185 185.680 ;
        RECT  0.600 183.850 64.400 185.680 ;
        RECT  46.230 183.720 51.730 185.870 ;
        RECT  54.855 183.850 56.700 185.950 ;
        RECT  4.895 155.120 7.525 171.290 ;
        RECT  8.170 155.125 8.490 171.290 ;
        RECT  22.160 155.160 22.510 171.290 ;
        RECT  22.810 155.140 23.130 171.290 ;
        RECT  49.615 155.125 51.855 171.290 ;
        RECT  52.795 155.295 53.105 171.290 ;
        RECT  53.655 155.035 53.935 171.290 ;
        RECT  56.365 155.280 56.645 171.315 ;
        RECT  57.120 155.300 57.400 171.315 ;
        RECT  57.835 155.130 58.115 171.315 ;
        RECT  0.600 155.310 64.400 171.290 ;
        RECT  56.240 155.310 61.880 171.315 ;
        RECT  53.895 155.310 55.870 171.370 ;
        RECT  3.220 155.310 3.500 171.380 ;
        RECT  34.655 155.310 38.715 171.480 ;
        RECT  39.605 155.310 42.020 171.480 ;
        RECT  2.000 0.000 63.000 60.210 ;
        RECT  0.600 0.600 64.400 60.210 ;
        RECT  0.600 0.600 1.210 135.520 ;
        RECT  0.600 91.020 64.400 135.520 ;
        RECT  4.080 91.020 60.940 135.690 ;
        RECT  62.580 91.020 62.995 135.710 ;
        LAYER M3 ;
        RECT  0.600 247.660 23.220 248.740 ;
        RECT  0.600 247.660 22.900 249.400 ;
        RECT  26.260 247.660 64.400 248.740 ;
        RECT  26.580 247.660 27.000 249.400 ;
        RECT  31.470 247.660 64.400 249.400 ;
        RECT  0.600 124.090 64.400 129.850 ;
        RECT  1.640 124.090 63.600 135.790 ;
        RECT  1.810 124.090 2.830 154.520 ;
        RECT  3.110 124.090 63.600 171.560 ;
        RECT  4.040 123.970 60.900 171.560 ;
        RECT  1.640 155.040 63.600 171.560 ;
        RECT  1.640 183.580 63.600 185.950 ;
        RECT  5.510 124.090 63.600 200.820 ;
        RECT  1.640 196.170 63.600 200.820 ;
        RECT  56.300 123.970 56.580 201.060 ;
        RECT  0.600 0.600 64.400 60.480 ;
        RECT  2.000 0.000 63.000 88.700 ;
        RECT  0.600 0.600 1.480 91.220 ;
        RECT  0.600 90.750 64.400 91.220 ;
        LAYER TOP_M ;
        RECT  0.600 247.690 64.400 248.850 ;
        RECT  0.600 247.690 23.010 249.400 ;
        RECT  26.470 247.690 27.110 249.400 ;
        RECT  31.360 247.690 64.400 249.400 ;
        RECT  2.000 0.000 63.000 91.190 ;
        RECT  0.600 0.600 64.400 91.190 ;
    END
END pc3b03d

MACRO pc3b03
    CLASS PAD ;
    FOREIGN pc3b03 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 65.000 BY 250.000 ;
    SYMMETRY X Y R90 ;
    SITE IOSite_c ;
    PIN PAD
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 55.440  LAYER TOP_M  ;
        ANTENNAPARTIALMETALSIDEAREA 287.938  LAYER M3  ;
        ANTENNAPARTIALMETALSIDEAREA 480.740  LAYER M2  ;
        ANTENNADIFFAREA 2657.280  LAYER TOP_M  ;
        ANTENNADIFFAREA 1209.600  LAYER M2  ;
        ANTENNADIFFAREA 2657.280  LAYER M3  ;
        ANTENNAPARTIALCUTAREA 632.318  LAYER TOP_V  ;
        ANTENNAPARTIALCUTAREA 349.898  LAYER V3  ;
        ANTENNAPARTIALCUTAREA 255.798  LAYER V2  ;
        PORT
        LAYER M3 ;
        RECT  23.740 249.580 25.740 250.000 ;
        LAYER M2 ;
        RECT  2.000 61.000 63.000 90.230 ;
        RECT  23.740 246.275 25.740 250.000 ;
        END
    END PAD
    PIN OEN
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 80.634  LAYER M2  ;
        ANTENNAPARTIALMETALSIDEAREA 41.679  LAYER M3  ;
        ANTENNAPARTIALMETALSIDEAREA 67.374  LAYER M1  ;
        ANTENNADIFFAREA 0.250  LAYER M3  ;
        ANTENNAPARTIALCUTAREA 0.203  LAYER V2  ;
        ANTENNAPARTIALCUTAREA 0.135  LAYER V3  ;
        ANTENNAGATEAREA 9.900  LAYER M3  ;
        ANTENNAGATEAREA 8.100  LAYER M2  ;
        PORT
        LAYER M3 ;
        RECT  29.900 249.580 30.630 250.000 ;
        LAYER M2 ;
        RECT  29.900 249.580 30.630 250.000 ;
        END
    END OEN
    PIN CIN
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 32.277  LAYER M3  ;
        ANTENNAPARTIALMETALSIDEAREA 96.916  LAYER M2  ;
        ANTENNAPARTIALMETALSIDEAREA 67.374  LAYER M1  ;
        ANTENNADIFFAREA 20.600  LAYER M3  ;
        ANTENNAPARTIALCUTAREA 0.135  LAYER V3  ;
        ANTENNAPARTIALCUTAREA 0.203  LAYER V2  ;
        PORT
        LAYER M3 ;
        RECT  28.870 249.580 29.600 250.000 ;
        LAYER M2 ;
        RECT  28.870 249.580 29.600 250.000 ;
        END
    END CIN
    PIN I
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 67.374  LAYER M1  ;
        ANTENNAPARTIALMETALSIDEAREA 80.804  LAYER M2  ;
        ANTENNAPARTIALMETALSIDEAREA 41.096  LAYER M3  ;
        ANTENNADIFFAREA 0.250  LAYER M3  ;
        ANTENNAPARTIALCUTAREA 0.270  LAYER V2  ;
        ANTENNAPARTIALCUTAREA 0.135  LAYER V3  ;
        ANTENNAGATEAREA 18.900  LAYER M2  ;
        ANTENNAGATEAREA 20.700  LAYER M3  ;
        PORT
        LAYER M3 ;
        RECT  27.840 249.580 28.570 250.000 ;
        LAYER M2 ;
        RECT  27.840 249.580 28.570 250.000 ;
        END
    END I
    PIN VDDO
        DIRECTION INOUT ;
        USE power ;
        PORT
        LAYER M3 ;
        RECT  64.200 192.330 65.000 200.640 ;
        RECT  0.000 201.660 65.000 221.520 ;
        RECT  0.000 222.720 65.000 246.820 ;
        RECT  0.000 192.330 0.800 200.640 ;
        LAYER M2 ;
        RECT  0.000 186.470 65.000 195.650 ;
        LAYER TOP_M ;
        RECT  0.000 195.170 65.000 200.640 ;
        RECT  0.000 201.660 65.000 221.520 ;
        RECT  0.000 222.720 65.000 246.820 ;
        END
    END VDDO
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        PORT
        LAYER M3 ;
        RECT  64.200 163.510 65.000 190.890 ;
        RECT  0.000 163.510 0.800 190.890 ;
        LAYER M2 ;
        RECT  0.000 172.080 65.000 183.060 ;
        LAYER TOP_M ;
        RECT  0.000 163.500 65.000 194.560 ;
        END
    END VDD
    PIN VSSO
        DIRECTION INOUT ;
        USE ground ;
        PORT
        LAYER M3 ;
        RECT  0.000 92.060 65.000 123.250 ;
        RECT  64.200 149.940 65.000 162.610 ;
        RECT  0.000 149.940 0.800 162.610 ;
        LAYER M2 ;
        RECT  0.000 147.040 65.000 154.520 ;
        LAYER TOP_M ;
        RECT  0.000 92.060 65.000 123.250 ;
        RECT  0.000 155.410 65.000 162.610 ;
        END
    END VSSO
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        PORT
        LAYER M3 ;
        RECT  64.200 130.690 65.000 148.880 ;
        RECT  0.000 130.690 0.800 148.880 ;
        LAYER M2 ;
        RECT  0.000 136.310 65.000 146.340 ;
        LAYER TOP_M ;
        RECT  0.000 123.850 65.000 154.560 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  2.000 0.000 63.000 250.000 ;
        RECT  0.000 88.990 65.000 130.360 ;
        RECT  0.000 136.510 65.000 157.550 ;
        RECT  0.315 158.150 64.700 158.460 ;
        RECT  0.300 158.930 64.700 159.230 ;
        RECT  0.300 159.530 64.700 159.830 ;
        RECT  0.300 160.130 64.700 160.430 ;
        RECT  0.300 160.730 64.700 161.030 ;
        RECT  0.300 161.330 64.700 161.630 ;
        RECT  0.300 161.910 64.700 162.190 ;
        RECT  0.300 162.490 64.700 162.770 ;
        RECT  0.300 163.070 64.700 163.350 ;
        RECT  0.300 163.650 64.700 163.950 ;
        RECT  0.300 164.250 64.700 164.550 ;
        RECT  0.300 164.850 64.700 165.150 ;
        RECT  0.300 165.450 64.700 165.750 ;
        RECT  0.300 166.050 64.700 166.350 ;
        RECT  0.300 166.650 64.700 166.960 ;
        RECT  0.300 167.260 64.700 167.560 ;
        RECT  0.300 167.860 64.700 168.160 ;
        RECT  0.000 169.150 65.000 197.240 ;
        RECT  0.600 0.600 64.400 250.000 ;
        RECT  0.000 198.470 65.000 250.000 ;
        LAYER M2 ;
        RECT  1.840 196.420 2.120 249.400 ;
        RECT  63.180 196.430 63.670 249.400 ;
        RECT  0.600 196.440 64.400 245.485 ;
        RECT  26.530 196.440 64.400 248.790 ;
        RECT  0.600 196.440 22.950 249.400 ;
        RECT  26.530 196.440 27.050 249.400 ;
        RECT  31.420 196.440 64.400 249.400 ;
        RECT  19.440 183.720 52.185 185.680 ;
        RECT  0.600 183.850 64.400 185.680 ;
        RECT  46.230 183.720 51.730 185.870 ;
        RECT  54.855 183.850 56.700 185.950 ;
        RECT  4.895 155.120 7.525 171.290 ;
        RECT  8.170 155.125 8.490 171.290 ;
        RECT  22.160 155.160 22.510 171.290 ;
        RECT  22.810 155.140 23.130 171.290 ;
        RECT  53.655 155.035 53.935 171.290 ;
        RECT  56.365 155.280 56.645 171.315 ;
        RECT  57.120 155.300 57.400 171.315 ;
        RECT  57.835 155.130 58.115 171.315 ;
        RECT  0.600 155.310 64.400 171.290 ;
        RECT  56.240 155.310 61.880 171.315 ;
        RECT  53.895 155.310 55.870 171.370 ;
        RECT  3.220 155.310 3.500 171.380 ;
        RECT  34.655 155.310 38.715 171.480 ;
        RECT  39.605 155.310 42.020 171.480 ;
        RECT  2.000 0.000 63.000 60.210 ;
        RECT  0.600 0.600 64.400 60.210 ;
        RECT  0.600 0.600 1.210 135.520 ;
        RECT  0.600 91.020 64.400 135.520 ;
        RECT  4.080 91.020 60.940 135.690 ;
        RECT  62.580 91.020 62.995 135.710 ;
        LAYER M3 ;
        RECT  0.600 247.660 23.220 248.740 ;
        RECT  0.600 247.660 22.900 249.400 ;
        RECT  26.260 247.660 64.400 248.740 ;
        RECT  26.580 247.660 27.000 249.400 ;
        RECT  31.470 247.660 64.400 249.400 ;
        RECT  0.600 124.090 64.400 129.850 ;
        RECT  1.640 124.090 63.600 135.790 ;
        RECT  1.810 124.090 2.830 154.520 ;
        RECT  3.110 124.090 63.600 171.560 ;
        RECT  4.040 123.970 60.900 171.560 ;
        RECT  1.640 155.040 63.600 171.560 ;
        RECT  1.640 183.580 63.600 185.950 ;
        RECT  5.510 124.090 63.600 200.820 ;
        RECT  1.640 196.170 63.600 200.820 ;
        RECT  56.300 123.970 56.580 201.060 ;
        RECT  0.600 0.600 64.400 60.480 ;
        RECT  2.000 0.000 63.000 88.700 ;
        RECT  0.600 0.600 1.480 91.220 ;
        RECT  0.600 90.750 64.400 91.220 ;
        LAYER TOP_M ;
        RECT  0.600 247.690 64.400 248.850 ;
        RECT  0.600 247.690 23.010 249.400 ;
        RECT  26.470 247.690 27.110 249.400 ;
        RECT  31.360 247.690 64.400 249.400 ;
        RECT  2.000 0.000 63.000 91.190 ;
        RECT  0.600 0.600 64.400 91.190 ;
    END
END pc3b03

MACRO pc3b02u
    CLASS PAD ;
    FOREIGN pc3b02u 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 65.000 BY 250.000 ;
    SYMMETRY X Y R90 ;
    SITE IOSite_c ;
    PIN PAD
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 55.440  LAYER TOP_M  ;
        ANTENNAPARTIALMETALSIDEAREA 287.938  LAYER M3  ;
        ANTENNAPARTIALMETALSIDEAREA 480.740  LAYER M2  ;
        ANTENNADIFFAREA 2657.280  LAYER TOP_M  ;
        ANTENNADIFFAREA 2657.280  LAYER M3  ;
        ANTENNADIFFAREA 1209.600  LAYER M2  ;
        ANTENNAPARTIALCUTAREA 632.318  LAYER TOP_V  ;
        ANTENNAPARTIALCUTAREA 349.898  LAYER V3  ;
        ANTENNAPARTIALCUTAREA 255.798  LAYER V2  ;
        PORT
        LAYER M3 ;
        RECT  23.740 249.580 25.740 250.000 ;
        LAYER M2 ;
        RECT  2.000 61.000 63.000 90.230 ;
        RECT  23.740 246.275 25.740 250.000 ;
        END
    END PAD
    PIN CIN
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 32.277  LAYER M3  ;
        ANTENNAPARTIALMETALSIDEAREA 96.916  LAYER M2  ;
        ANTENNAPARTIALMETALSIDEAREA 67.374  LAYER M1  ;
        ANTENNADIFFAREA 20.600  LAYER M3  ;
        ANTENNAPARTIALCUTAREA 0.135  LAYER V3  ;
        ANTENNAPARTIALCUTAREA 0.203  LAYER V2  ;
        PORT
        LAYER M3 ;
        RECT  28.870 249.580 29.600 250.000 ;
        LAYER M2 ;
        RECT  28.870 249.580 29.600 250.000 ;
        END
    END CIN
    PIN OEN
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 80.634  LAYER M2  ;
        ANTENNAPARTIALMETALSIDEAREA 67.374  LAYER M1  ;
        ANTENNAPARTIALMETALSIDEAREA 41.679  LAYER M3  ;
        ANTENNADIFFAREA 0.250  LAYER M3  ;
        ANTENNAPARTIALCUTAREA 0.203  LAYER V2  ;
        ANTENNAPARTIALCUTAREA 0.135  LAYER V3  ;
        ANTENNAGATEAREA 8.100  LAYER M2  ;
        ANTENNAGATEAREA 9.900  LAYER M3  ;
        PORT
        LAYER M3 ;
        RECT  29.900 249.580 30.630 250.000 ;
        LAYER M2 ;
        RECT  29.900 249.580 30.630 250.000 ;
        END
    END OEN
    PIN I
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 67.374  LAYER M1  ;
        ANTENNAPARTIALMETALSIDEAREA 80.804  LAYER M2  ;
        ANTENNAPARTIALMETALSIDEAREA 41.096  LAYER M3  ;
        ANTENNADIFFAREA 0.250  LAYER M3  ;
        ANTENNAPARTIALCUTAREA 0.270  LAYER V2  ;
        ANTENNAPARTIALCUTAREA 0.135  LAYER V3  ;
        ANTENNAGATEAREA 18.900  LAYER M2  ;
        ANTENNAGATEAREA 20.700  LAYER M3  ;
        PORT
        LAYER M3 ;
        RECT  27.840 249.580 28.570 250.000 ;
        LAYER M2 ;
        RECT  27.840 249.580 28.570 250.000 ;
        END
    END I
    PIN VDDO
        DIRECTION INOUT ;
        USE power ;
        PORT
        LAYER M3 ;
        RECT  64.200 192.330 65.000 200.640 ;
        RECT  0.000 201.660 65.000 221.520 ;
        RECT  0.000 222.720 65.000 246.820 ;
        RECT  0.000 192.330 0.800 200.640 ;
        LAYER M2 ;
        RECT  0.000 186.470 65.000 195.650 ;
        LAYER TOP_M ;
        RECT  0.000 195.170 65.000 200.640 ;
        RECT  0.000 201.660 65.000 221.520 ;
        RECT  0.000 222.720 65.000 246.820 ;
        END
    END VDDO
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        PORT
        LAYER M3 ;
        RECT  64.200 163.510 65.000 190.890 ;
        RECT  0.000 163.510 0.800 190.890 ;
        LAYER M2 ;
        RECT  0.000 172.080 65.000 183.060 ;
        LAYER TOP_M ;
        RECT  0.000 163.500 65.000 194.560 ;
        END
    END VDD
    PIN VSSO
        DIRECTION INOUT ;
        USE ground ;
        PORT
        LAYER M3 ;
        RECT  0.000 92.060 65.000 123.250 ;
        RECT  64.200 149.940 65.000 162.610 ;
        RECT  0.000 149.940 0.800 162.610 ;
        LAYER M2 ;
        RECT  0.000 147.040 65.000 154.520 ;
        LAYER TOP_M ;
        RECT  0.000 92.060 65.000 123.250 ;
        RECT  0.000 155.410 65.000 162.610 ;
        END
    END VSSO
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        PORT
        LAYER M3 ;
        RECT  64.200 130.690 65.000 148.880 ;
        RECT  0.000 130.690 0.800 148.880 ;
        LAYER M2 ;
        RECT  0.000 136.310 65.000 146.340 ;
        LAYER TOP_M ;
        RECT  0.000 123.850 65.000 154.560 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  2.000 0.000 63.000 250.000 ;
        RECT  0.000 88.990 65.000 130.360 ;
        RECT  0.000 136.510 65.000 157.550 ;
        RECT  0.315 158.150 64.700 158.460 ;
        RECT  0.300 158.930 64.700 159.230 ;
        RECT  0.300 159.530 64.700 159.830 ;
        RECT  0.300 160.130 64.700 160.430 ;
        RECT  0.300 160.730 64.700 161.030 ;
        RECT  0.300 161.330 64.700 161.630 ;
        RECT  0.300 161.910 64.700 162.190 ;
        RECT  0.300 162.490 64.700 162.770 ;
        RECT  0.300 163.070 64.700 163.350 ;
        RECT  0.300 163.650 64.700 163.950 ;
        RECT  0.300 164.250 64.700 164.550 ;
        RECT  0.300 164.850 64.700 165.150 ;
        RECT  0.300 165.450 64.700 165.750 ;
        RECT  0.300 166.050 64.700 166.350 ;
        RECT  0.300 166.650 64.700 166.960 ;
        RECT  0.300 167.260 64.700 167.560 ;
        RECT  0.300 167.860 64.700 168.160 ;
        RECT  0.000 169.150 65.000 197.240 ;
        RECT  0.600 0.600 64.400 250.000 ;
        RECT  0.000 198.470 65.000 250.000 ;
        LAYER M2 ;
        RECT  1.840 196.420 2.120 249.400 ;
        RECT  63.180 196.430 63.670 249.400 ;
        RECT  0.600 196.440 64.400 245.485 ;
        RECT  26.530 196.440 64.400 248.790 ;
        RECT  0.600 196.440 22.950 249.400 ;
        RECT  26.530 196.440 27.050 249.400 ;
        RECT  31.420 196.440 64.400 249.400 ;
        RECT  18.205 183.720 52.025 185.680 ;
        RECT  0.600 183.850 64.400 185.680 ;
        RECT  46.230 183.720 51.730 185.870 ;
        RECT  54.940 183.850 56.670 185.870 ;
        RECT  8.735 155.125 9.055 171.290 ;
        RECT  21.065 155.160 21.415 171.290 ;
        RECT  21.715 155.140 22.035 171.290 ;
        RECT  53.655 155.035 53.935 171.290 ;
        RECT  56.365 155.280 56.645 171.315 ;
        RECT  57.120 155.300 57.400 171.315 ;
        RECT  57.835 155.130 58.115 171.315 ;
        RECT  0.600 155.310 64.400 171.290 ;
        RECT  56.240 155.310 61.880 171.315 ;
        RECT  53.895 155.310 55.870 171.370 ;
        RECT  32.965 155.310 33.465 171.375 ;
        RECT  3.220 155.310 3.500 171.380 ;
        RECT  34.655 155.310 38.715 171.480 ;
        RECT  39.605 155.310 42.020 171.480 ;
        RECT  2.000 0.000 63.000 60.210 ;
        RECT  0.600 0.600 64.400 60.210 ;
        RECT  0.600 0.600 1.210 135.520 ;
        RECT  0.600 91.020 64.400 135.520 ;
        RECT  4.080 91.020 60.940 135.690 ;
        RECT  62.580 91.020 62.995 135.710 ;
        LAYER M3 ;
        RECT  0.600 247.660 23.220 248.740 ;
        RECT  0.600 247.660 22.900 249.400 ;
        RECT  26.260 247.660 64.400 248.740 ;
        RECT  26.580 247.660 27.000 249.400 ;
        RECT  31.470 247.660 64.400 249.400 ;
        RECT  0.600 124.090 64.400 129.850 ;
        RECT  1.640 124.090 63.600 135.790 ;
        RECT  1.810 124.090 2.830 154.520 ;
        RECT  3.110 124.090 63.600 171.560 ;
        RECT  4.040 123.970 60.900 171.560 ;
        RECT  1.640 155.040 63.600 171.560 ;
        RECT  1.640 183.580 63.600 185.950 ;
        RECT  5.490 124.090 63.600 200.820 ;
        RECT  1.640 196.170 63.600 200.820 ;
        RECT  56.300 123.970 56.580 201.060 ;
        RECT  0.600 0.600 64.400 60.480 ;
        RECT  2.000 0.000 63.000 88.700 ;
        RECT  0.600 0.600 1.480 91.220 ;
        RECT  0.600 90.750 64.400 91.220 ;
        LAYER TOP_M ;
        RECT  0.600 247.690 64.400 248.850 ;
        RECT  0.600 247.690 23.010 249.400 ;
        RECT  26.470 247.690 27.110 249.400 ;
        RECT  31.360 247.690 64.400 249.400 ;
        RECT  2.000 0.000 63.000 91.190 ;
        RECT  0.600 0.600 64.400 91.190 ;
    END
END pc3b02u

MACRO pc3b02d
    CLASS PAD ;
    FOREIGN pc3b02d 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 65.000 BY 250.000 ;
    SYMMETRY X Y R90 ;
    SITE IOSite_c ;
    PIN PAD
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 55.440  LAYER TOP_M  ;
        ANTENNAPARTIALMETALSIDEAREA 287.938  LAYER M3  ;
        ANTENNAPARTIALMETALSIDEAREA 480.740  LAYER M2  ;
        ANTENNADIFFAREA 2657.280  LAYER TOP_M  ;
        ANTENNADIFFAREA 2657.280  LAYER M3  ;
        ANTENNADIFFAREA 1209.600  LAYER M2  ;
        ANTENNAPARTIALCUTAREA 632.318  LAYER TOP_V  ;
        ANTENNAPARTIALCUTAREA 349.898  LAYER V3  ;
        ANTENNAPARTIALCUTAREA 255.798  LAYER V2  ;
        PORT
        LAYER M3 ;
        RECT  23.740 249.580 25.740 250.000 ;
        LAYER M2 ;
        RECT  2.000 61.000 63.000 90.230 ;
        RECT  23.740 246.275 25.740 250.000 ;
        END
    END PAD
    PIN CIN
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 32.277  LAYER M3  ;
        ANTENNAPARTIALMETALSIDEAREA 96.916  LAYER M2  ;
        ANTENNAPARTIALMETALSIDEAREA 67.374  LAYER M1  ;
        ANTENNADIFFAREA 20.600  LAYER M3  ;
        ANTENNAPARTIALCUTAREA 0.135  LAYER V3  ;
        ANTENNAPARTIALCUTAREA 0.203  LAYER V2  ;
        PORT
        LAYER M3 ;
        RECT  28.870 249.580 29.600 250.000 ;
        LAYER M2 ;
        RECT  28.870 249.580 29.600 250.000 ;
        END
    END CIN
    PIN OEN
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 80.634  LAYER M2  ;
        ANTENNAPARTIALMETALSIDEAREA 67.374  LAYER M1  ;
        ANTENNAPARTIALMETALSIDEAREA 41.679  LAYER M3  ;
        ANTENNADIFFAREA 0.250  LAYER M3  ;
        ANTENNAPARTIALCUTAREA 0.203  LAYER V2  ;
        ANTENNAPARTIALCUTAREA 0.135  LAYER V3  ;
        ANTENNAGATEAREA 8.100  LAYER M2  ;
        ANTENNAGATEAREA 9.900  LAYER M3  ;
        PORT
        LAYER M3 ;
        RECT  29.900 249.580 30.630 250.000 ;
        LAYER M2 ;
        RECT  29.900 249.580 30.630 250.000 ;
        END
    END OEN
    PIN I
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 67.374  LAYER M1  ;
        ANTENNAPARTIALMETALSIDEAREA 80.804  LAYER M2  ;
        ANTENNAPARTIALMETALSIDEAREA 41.096  LAYER M3  ;
        ANTENNADIFFAREA 0.250  LAYER M3  ;
        ANTENNAPARTIALCUTAREA 0.270  LAYER V2  ;
        ANTENNAPARTIALCUTAREA 0.135  LAYER V3  ;
        ANTENNAGATEAREA 18.900  LAYER M2  ;
        ANTENNAGATEAREA 20.700  LAYER M3  ;
        PORT
        LAYER M3 ;
        RECT  27.840 249.580 28.570 250.000 ;
        LAYER M2 ;
        RECT  27.840 249.580 28.570 250.000 ;
        END
    END I
    PIN VDDO
        DIRECTION INOUT ;
        USE power ;
        PORT
        LAYER M3 ;
        RECT  64.200 192.330 65.000 200.640 ;
        RECT  0.000 201.660 65.000 221.520 ;
        RECT  0.000 222.720 65.000 246.820 ;
        RECT  0.000 192.330 0.800 200.640 ;
        LAYER M2 ;
        RECT  0.000 186.470 65.000 195.650 ;
        LAYER TOP_M ;
        RECT  0.000 195.170 65.000 200.640 ;
        RECT  0.000 201.660 65.000 221.520 ;
        RECT  0.000 222.720 65.000 246.820 ;
        END
    END VDDO
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        PORT
        LAYER M3 ;
        RECT  64.200 163.510 65.000 190.890 ;
        RECT  0.000 163.510 0.800 190.890 ;
        LAYER M2 ;
        RECT  0.000 172.080 65.000 183.060 ;
        LAYER TOP_M ;
        RECT  0.000 163.500 65.000 194.560 ;
        END
    END VDD
    PIN VSSO
        DIRECTION INOUT ;
        USE ground ;
        PORT
        LAYER M3 ;
        RECT  0.000 92.060 65.000 123.250 ;
        RECT  64.200 149.940 65.000 162.610 ;
        RECT  0.000 149.940 0.800 162.610 ;
        LAYER M2 ;
        RECT  0.000 147.040 65.000 154.520 ;
        LAYER TOP_M ;
        RECT  0.000 92.060 65.000 123.250 ;
        RECT  0.000 155.410 65.000 162.610 ;
        END
    END VSSO
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        PORT
        LAYER M3 ;
        RECT  64.200 130.690 65.000 148.880 ;
        RECT  0.000 130.690 0.800 148.880 ;
        LAYER M2 ;
        RECT  0.000 136.310 65.000 146.340 ;
        LAYER TOP_M ;
        RECT  0.000 123.850 65.000 154.560 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  2.000 0.000 63.000 250.000 ;
        RECT  0.000 88.990 65.000 130.360 ;
        RECT  0.000 136.510 65.000 157.550 ;
        RECT  0.315 158.150 64.700 158.460 ;
        RECT  0.300 158.930 64.700 159.230 ;
        RECT  0.300 159.530 64.700 159.830 ;
        RECT  0.300 160.130 64.700 160.430 ;
        RECT  0.300 160.730 64.700 161.030 ;
        RECT  0.300 161.330 64.700 161.630 ;
        RECT  0.300 161.910 64.700 162.190 ;
        RECT  0.300 162.490 64.700 162.770 ;
        RECT  0.300 163.070 64.700 163.350 ;
        RECT  0.300 163.650 64.700 163.950 ;
        RECT  0.300 164.250 64.700 164.550 ;
        RECT  0.300 164.850 64.700 165.150 ;
        RECT  0.300 165.450 64.700 165.750 ;
        RECT  0.300 166.050 64.700 166.350 ;
        RECT  0.300 166.650 64.700 166.960 ;
        RECT  0.300 167.260 64.700 167.560 ;
        RECT  0.300 167.860 64.700 168.160 ;
        RECT  0.000 169.150 65.000 197.240 ;
        RECT  0.600 0.600 64.400 250.000 ;
        RECT  0.000 198.470 65.000 250.000 ;
        LAYER M2 ;
        RECT  1.840 196.420 2.120 249.400 ;
        RECT  63.180 196.430 63.670 249.400 ;
        RECT  0.600 196.440 64.400 245.485 ;
        RECT  26.530 196.440 64.400 248.790 ;
        RECT  0.600 196.440 22.950 249.400 ;
        RECT  26.530 196.440 27.050 249.400 ;
        RECT  31.420 196.440 64.400 249.400 ;
        RECT  18.205 183.720 52.025 185.680 ;
        RECT  0.600 183.850 64.400 185.680 ;
        RECT  46.230 183.720 51.730 185.870 ;
        RECT  54.940 183.850 56.670 185.870 ;
        RECT  8.735 155.125 9.055 171.290 ;
        RECT  21.065 155.160 21.415 171.290 ;
        RECT  21.715 155.140 22.035 171.290 ;
        RECT  49.535 155.125 51.775 171.290 ;
        RECT  52.715 155.295 53.025 171.290 ;
        RECT  53.655 155.035 53.935 171.290 ;
        RECT  56.365 155.280 56.645 171.315 ;
        RECT  57.120 155.300 57.400 171.315 ;
        RECT  57.835 155.130 58.115 171.315 ;
        RECT  0.600 155.310 64.400 171.290 ;
        RECT  56.240 155.310 61.880 171.315 ;
        RECT  53.895 155.310 55.870 171.370 ;
        RECT  3.220 155.310 3.500 171.380 ;
        RECT  34.655 155.310 38.715 171.480 ;
        RECT  39.605 155.310 42.020 171.480 ;
        RECT  2.000 0.000 63.000 60.210 ;
        RECT  0.600 0.600 64.400 60.210 ;
        RECT  0.600 0.600 1.210 135.520 ;
        RECT  0.600 91.020 64.400 135.520 ;
        RECT  4.080 91.020 60.940 135.690 ;
        RECT  62.580 91.020 62.995 135.710 ;
        LAYER M3 ;
        RECT  0.600 247.660 23.220 248.740 ;
        RECT  0.600 247.660 22.900 249.400 ;
        RECT  26.260 247.660 64.400 248.740 ;
        RECT  26.580 247.660 27.000 249.400 ;
        RECT  31.470 247.660 64.400 249.400 ;
        RECT  0.600 124.090 64.400 129.850 ;
        RECT  1.640 124.090 63.600 135.790 ;
        RECT  1.810 124.090 2.830 154.520 ;
        RECT  3.110 124.090 63.600 171.560 ;
        RECT  4.040 123.970 60.900 171.560 ;
        RECT  1.640 155.040 63.600 171.560 ;
        RECT  1.640 183.580 63.600 185.950 ;
        RECT  5.490 124.090 63.600 200.820 ;
        RECT  1.640 196.170 63.600 200.820 ;
        RECT  56.300 123.970 56.580 201.060 ;
        RECT  0.600 0.600 64.400 60.480 ;
        RECT  2.000 0.000 63.000 88.700 ;
        RECT  0.600 0.600 1.480 91.220 ;
        RECT  0.600 90.750 64.400 91.220 ;
        LAYER TOP_M ;
        RECT  0.600 247.690 64.400 248.850 ;
        RECT  0.600 247.690 23.010 249.400 ;
        RECT  26.470 247.690 27.110 249.400 ;
        RECT  31.360 247.690 64.400 249.400 ;
        RECT  2.000 0.000 63.000 91.190 ;
        RECT  0.600 0.600 64.400 91.190 ;
    END
END pc3b02d

MACRO pc3b02
    CLASS PAD ;
    FOREIGN pc3b02 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 65.000 BY 250.000 ;
    SYMMETRY X Y R90 ;
    SITE IOSite_c ;
    PIN PAD
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 55.440  LAYER TOP_M  ;
        ANTENNAPARTIALMETALSIDEAREA 287.938  LAYER M3  ;
        ANTENNAPARTIALMETALSIDEAREA 480.740  LAYER M2  ;
        ANTENNADIFFAREA 2657.280  LAYER TOP_M  ;
        ANTENNADIFFAREA 2657.280  LAYER M3  ;
        ANTENNADIFFAREA 1209.600  LAYER M2  ;
        ANTENNAPARTIALCUTAREA 632.318  LAYER TOP_V  ;
        ANTENNAPARTIALCUTAREA 349.898  LAYER V3  ;
        ANTENNAPARTIALCUTAREA 255.798  LAYER V2  ;
        PORT
        LAYER M3 ;
        RECT  23.740 249.580 25.740 250.000 ;
        LAYER M2 ;
        RECT  2.000 61.000 63.000 90.230 ;
        RECT  23.740 246.275 25.740 250.000 ;
        END
    END PAD
    PIN CIN
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 32.277  LAYER M3  ;
        ANTENNAPARTIALMETALSIDEAREA 96.916  LAYER M2  ;
        ANTENNAPARTIALMETALSIDEAREA 67.374  LAYER M1  ;
        ANTENNADIFFAREA 20.600  LAYER M3  ;
        ANTENNAPARTIALCUTAREA 0.135  LAYER V3  ;
        ANTENNAPARTIALCUTAREA 0.203  LAYER V2  ;
        PORT
        LAYER M3 ;
        RECT  28.870 249.580 29.600 250.000 ;
        LAYER M2 ;
        RECT  28.870 249.580 29.600 250.000 ;
        END
    END CIN
    PIN OEN
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 80.634  LAYER M2  ;
        ANTENNAPARTIALMETALSIDEAREA 67.374  LAYER M1  ;
        ANTENNAPARTIALMETALSIDEAREA 41.679  LAYER M3  ;
        ANTENNADIFFAREA 0.250  LAYER M3  ;
        ANTENNAPARTIALCUTAREA 0.203  LAYER V2  ;
        ANTENNAPARTIALCUTAREA 0.135  LAYER V3  ;
        ANTENNAGATEAREA 8.100  LAYER M2  ;
        ANTENNAGATEAREA 9.900  LAYER M3  ;
        PORT
        LAYER M3 ;
        RECT  29.900 249.580 30.630 250.000 ;
        LAYER M2 ;
        RECT  29.900 249.580 30.630 250.000 ;
        END
    END OEN
    PIN I
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 67.374  LAYER M1  ;
        ANTENNAPARTIALMETALSIDEAREA 80.804  LAYER M2  ;
        ANTENNAPARTIALMETALSIDEAREA 41.096  LAYER M3  ;
        ANTENNADIFFAREA 0.250  LAYER M3  ;
        ANTENNAPARTIALCUTAREA 0.270  LAYER V2  ;
        ANTENNAPARTIALCUTAREA 0.135  LAYER V3  ;
        ANTENNAGATEAREA 18.900  LAYER M2  ;
        ANTENNAGATEAREA 20.700  LAYER M3  ;
        PORT
        LAYER M3 ;
        RECT  27.840 249.580 28.570 250.000 ;
        LAYER M2 ;
        RECT  27.840 249.580 28.570 250.000 ;
        END
    END I
    PIN VDDO
        DIRECTION INOUT ;
        USE power ;
        PORT
        LAYER M3 ;
        RECT  64.200 192.330 65.000 200.640 ;
        RECT  0.000 201.660 65.000 221.520 ;
        RECT  0.000 222.720 65.000 246.820 ;
        RECT  0.000 192.330 0.800 200.640 ;
        LAYER M2 ;
        RECT  0.000 186.470 65.000 195.650 ;
        LAYER TOP_M ;
        RECT  0.000 195.170 65.000 200.640 ;
        RECT  0.000 201.660 65.000 221.520 ;
        RECT  0.000 222.720 65.000 246.820 ;
        END
    END VDDO
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        PORT
        LAYER M3 ;
        RECT  64.200 163.510 65.000 190.890 ;
        RECT  0.000 163.510 0.800 190.890 ;
        LAYER M2 ;
        RECT  0.000 172.080 65.000 183.060 ;
        LAYER TOP_M ;
        RECT  0.000 163.500 65.000 194.560 ;
        END
    END VDD
    PIN VSSO
        DIRECTION INOUT ;
        USE ground ;
        PORT
        LAYER M3 ;
        RECT  0.000 92.060 65.000 123.250 ;
        RECT  64.200 149.940 65.000 162.610 ;
        RECT  0.000 149.940 0.800 162.610 ;
        LAYER M2 ;
        RECT  0.000 147.040 65.000 154.520 ;
        LAYER TOP_M ;
        RECT  0.000 92.060 65.000 123.250 ;
        RECT  0.000 155.410 65.000 162.610 ;
        END
    END VSSO
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        PORT
        LAYER M3 ;
        RECT  64.200 130.690 65.000 148.880 ;
        RECT  0.000 130.690 0.800 148.880 ;
        LAYER M2 ;
        RECT  0.000 136.310 65.000 146.340 ;
        LAYER TOP_M ;
        RECT  0.000 123.850 65.000 154.560 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  2.000 0.000 63.000 250.000 ;
        RECT  0.000 88.990 65.000 130.360 ;
        RECT  0.000 136.510 65.000 157.550 ;
        RECT  0.315 158.150 64.700 158.460 ;
        RECT  0.300 158.930 64.700 159.230 ;
        RECT  0.300 159.530 64.700 159.830 ;
        RECT  0.300 160.130 64.700 160.430 ;
        RECT  0.300 160.730 64.700 161.030 ;
        RECT  0.300 161.330 64.700 161.630 ;
        RECT  0.300 161.910 64.700 162.190 ;
        RECT  0.300 162.490 64.700 162.770 ;
        RECT  0.300 163.070 64.700 163.350 ;
        RECT  0.300 163.650 64.700 163.950 ;
        RECT  0.300 164.250 64.700 164.550 ;
        RECT  0.300 164.850 64.700 165.150 ;
        RECT  0.300 165.450 64.700 165.750 ;
        RECT  0.300 166.050 64.700 166.350 ;
        RECT  0.300 166.650 64.700 166.960 ;
        RECT  0.300 167.260 64.700 167.560 ;
        RECT  0.300 167.860 64.700 168.160 ;
        RECT  0.000 169.150 65.000 197.240 ;
        RECT  0.600 0.600 64.400 250.000 ;
        RECT  0.000 198.470 65.000 250.000 ;
        LAYER M2 ;
        RECT  1.840 196.420 2.120 249.400 ;
        RECT  63.180 196.430 63.670 249.400 ;
        RECT  0.600 196.440 64.400 245.485 ;
        RECT  26.530 196.440 64.400 248.790 ;
        RECT  0.600 196.440 22.950 249.400 ;
        RECT  26.530 196.440 27.050 249.400 ;
        RECT  31.420 196.440 64.400 249.400 ;
        RECT  18.205 183.720 52.025 185.680 ;
        RECT  0.600 183.850 64.400 185.680 ;
        RECT  46.230 183.720 51.730 185.870 ;
        RECT  54.940 183.850 56.670 185.870 ;
        RECT  8.735 155.125 9.055 171.290 ;
        RECT  21.065 155.160 21.415 171.290 ;
        RECT  21.715 155.140 22.035 171.290 ;
        RECT  53.655 155.035 53.935 171.290 ;
        RECT  56.365 155.280 56.645 171.315 ;
        RECT  57.120 155.300 57.400 171.315 ;
        RECT  57.835 155.130 58.115 171.315 ;
        RECT  0.600 155.310 64.400 171.290 ;
        RECT  56.240 155.310 61.880 171.315 ;
        RECT  53.895 155.310 55.870 171.370 ;
        RECT  3.220 155.310 3.500 171.380 ;
        RECT  34.655 155.310 38.715 171.480 ;
        RECT  39.605 155.310 42.020 171.480 ;
        RECT  2.000 0.000 63.000 60.210 ;
        RECT  0.600 0.600 64.400 60.210 ;
        RECT  0.600 0.600 1.210 135.520 ;
        RECT  0.600 91.020 64.400 135.520 ;
        RECT  4.080 91.020 60.940 135.690 ;
        RECT  62.580 91.020 62.995 135.710 ;
        LAYER M3 ;
        RECT  0.600 247.660 23.220 248.740 ;
        RECT  0.600 247.660 22.900 249.400 ;
        RECT  26.260 247.660 64.400 248.740 ;
        RECT  26.580 247.660 27.000 249.400 ;
        RECT  31.470 247.660 64.400 249.400 ;
        RECT  0.600 124.090 64.400 129.850 ;
        RECT  1.640 124.090 63.600 135.790 ;
        RECT  1.810 124.090 2.830 154.520 ;
        RECT  3.110 124.090 63.600 171.560 ;
        RECT  4.040 123.970 60.900 171.560 ;
        RECT  1.640 155.040 63.600 171.560 ;
        RECT  1.640 183.580 63.600 185.950 ;
        RECT  5.490 124.090 63.600 200.820 ;
        RECT  1.640 196.170 63.600 200.820 ;
        RECT  56.300 123.970 56.580 201.060 ;
        RECT  0.600 0.600 64.400 60.480 ;
        RECT  2.000 0.000 63.000 88.700 ;
        RECT  0.600 0.600 1.480 91.220 ;
        RECT  0.600 90.750 64.400 91.220 ;
        LAYER TOP_M ;
        RECT  0.600 247.690 64.400 248.850 ;
        RECT  0.600 247.690 23.010 249.400 ;
        RECT  26.470 247.690 27.110 249.400 ;
        RECT  31.360 247.690 64.400 249.400 ;
        RECT  2.000 0.000 63.000 91.190 ;
        RECT  0.600 0.600 64.400 91.190 ;
    END
END pc3b02

MACRO pc3b01u
    CLASS PAD ;
    FOREIGN pc3b01u 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 65.000 BY 250.000 ;
    SYMMETRY X Y R90 ;
    SITE IOSite_c ;
    PIN PAD
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 55.440  LAYER TOP_M  ;
        ANTENNAPARTIALMETALSIDEAREA 287.938  LAYER M3  ;
        ANTENNAPARTIALMETALSIDEAREA 480.740  LAYER M2  ;
        ANTENNADIFFAREA 2657.280  LAYER TOP_M  ;
        ANTENNADIFFAREA 2657.280  LAYER M3  ;
        ANTENNADIFFAREA 1209.600  LAYER M2  ;
        ANTENNAPARTIALCUTAREA 632.318  LAYER TOP_V  ;
        ANTENNAPARTIALCUTAREA 349.898  LAYER V3  ;
        ANTENNAPARTIALCUTAREA 255.798  LAYER V2  ;
        PORT
        LAYER M3 ;
        RECT  23.740 249.580 25.740 250.000 ;
        LAYER M2 ;
        RECT  2.000 61.000 63.000 90.230 ;
        RECT  23.740 246.275 25.740 250.000 ;
        END
    END PAD
    PIN OEN
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 67.374  LAYER M1  ;
        ANTENNAPARTIALMETALSIDEAREA 80.634  LAYER M2  ;
        ANTENNAPARTIALMETALSIDEAREA 41.679  LAYER M3  ;
        ANTENNADIFFAREA 0.250  LAYER M3  ;
        ANTENNAPARTIALCUTAREA 0.203  LAYER V2  ;
        ANTENNAPARTIALCUTAREA 0.135  LAYER V3  ;
        ANTENNAGATEAREA 8.100  LAYER M2  ;
        ANTENNAGATEAREA 9.900  LAYER M3  ;
        PORT
        LAYER M3 ;
        RECT  29.900 249.580 30.630 250.000 ;
        LAYER M2 ;
        RECT  29.900 249.580 30.630 250.000 ;
        END
    END OEN
    PIN CIN
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 32.277  LAYER M3  ;
        ANTENNAPARTIALMETALSIDEAREA 96.916  LAYER M2  ;
        ANTENNAPARTIALMETALSIDEAREA 67.374  LAYER M1  ;
        ANTENNADIFFAREA 20.600  LAYER M3  ;
        ANTENNAPARTIALCUTAREA 0.135  LAYER V3  ;
        ANTENNAPARTIALCUTAREA 0.203  LAYER V2  ;
        PORT
        LAYER M3 ;
        RECT  28.870 249.580 29.600 250.000 ;
        LAYER M2 ;
        RECT  28.870 249.580 29.600 250.000 ;
        END
    END CIN
    PIN I
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 80.804  LAYER M2  ;
        ANTENNAPARTIALMETALSIDEAREA 67.374  LAYER M1  ;
        ANTENNAPARTIALMETALSIDEAREA 41.096  LAYER M3  ;
        ANTENNADIFFAREA 0.250  LAYER M3  ;
        ANTENNAPARTIALCUTAREA 0.203  LAYER V2  ;
        ANTENNAPARTIALCUTAREA 0.135  LAYER V3  ;
        ANTENNAGATEAREA 8.100  LAYER M2  ;
        ANTENNAGATEAREA 9.900  LAYER M3  ;
        PORT
        LAYER M3 ;
        RECT  27.840 249.580 28.570 250.000 ;
        LAYER M2 ;
        RECT  27.840 249.580 28.570 250.000 ;
        END
    END I
    PIN VDDO
        DIRECTION INOUT ;
        USE power ;
        PORT
        LAYER M3 ;
        RECT  64.200 192.330 65.000 200.640 ;
        RECT  0.000 201.660 65.000 221.520 ;
        RECT  0.000 222.720 65.000 246.820 ;
        RECT  0.000 192.330 0.800 200.640 ;
        LAYER M2 ;
        RECT  0.000 186.470 65.000 195.650 ;
        LAYER TOP_M ;
        RECT  0.000 195.170 65.000 200.640 ;
        RECT  0.000 201.660 65.000 221.520 ;
        RECT  0.000 222.720 65.000 246.820 ;
        END
    END VDDO
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        PORT
        LAYER M3 ;
        RECT  64.200 163.510 65.000 190.890 ;
        RECT  0.000 163.510 0.800 190.890 ;
        LAYER M2 ;
        RECT  0.000 172.080 65.000 183.060 ;
        LAYER TOP_M ;
        RECT  0.000 163.500 65.000 194.560 ;
        END
    END VDD
    PIN VSSO
        DIRECTION INOUT ;
        USE ground ;
        PORT
        LAYER M3 ;
        RECT  0.000 92.060 65.000 123.250 ;
        RECT  64.200 149.940 65.000 162.610 ;
        RECT  0.000 149.940 0.800 162.610 ;
        LAYER M2 ;
        RECT  0.000 147.040 65.000 154.520 ;
        LAYER TOP_M ;
        RECT  0.000 92.060 65.000 123.250 ;
        RECT  0.000 155.410 65.000 162.610 ;
        END
    END VSSO
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        PORT
        LAYER M3 ;
        RECT  64.200 130.690 65.000 148.880 ;
        RECT  0.000 130.690 0.800 148.880 ;
        LAYER M2 ;
        RECT  0.000 136.310 65.000 146.340 ;
        LAYER TOP_M ;
        RECT  0.000 123.850 65.000 154.560 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  2.000 0.000 63.000 250.000 ;
        RECT  0.000 88.990 65.000 130.360 ;
        RECT  0.000 136.510 65.000 157.550 ;
        RECT  0.315 158.150 64.700 158.460 ;
        RECT  0.300 158.930 64.700 159.230 ;
        RECT  0.300 159.530 64.700 159.830 ;
        RECT  0.300 160.130 64.700 160.430 ;
        RECT  0.300 160.730 64.700 161.030 ;
        RECT  0.300 161.330 64.700 161.630 ;
        RECT  0.300 161.910 64.700 162.190 ;
        RECT  0.300 162.490 64.700 162.770 ;
        RECT  0.300 163.070 64.700 163.350 ;
        RECT  0.300 163.650 64.700 163.950 ;
        RECT  0.300 164.250 64.700 164.550 ;
        RECT  0.300 164.850 64.700 165.150 ;
        RECT  0.300 165.450 64.700 165.750 ;
        RECT  0.300 166.050 64.700 166.350 ;
        RECT  0.300 166.650 64.700 166.960 ;
        RECT  0.300 167.260 64.700 167.560 ;
        RECT  0.300 167.860 64.700 168.160 ;
        RECT  0.000 169.150 65.000 197.240 ;
        RECT  0.600 0.600 64.400 250.000 ;
        RECT  0.000 198.470 65.000 250.000 ;
        LAYER M2 ;
        RECT  1.840 196.420 2.120 249.400 ;
        RECT  63.180 196.430 63.670 249.400 ;
        RECT  0.600 196.440 64.400 245.485 ;
        RECT  26.530 196.440 64.400 248.790 ;
        RECT  0.600 196.440 22.950 249.400 ;
        RECT  26.530 196.440 27.050 249.400 ;
        RECT  31.420 196.440 64.400 249.400 ;
        RECT  14.290 183.720 52.380 185.680 ;
        RECT  0.600 183.850 64.400 185.680 ;
        RECT  54.910 183.850 57.160 185.865 ;
        RECT  46.230 183.720 51.730 185.870 ;
        RECT  18.450 155.160 18.800 171.290 ;
        RECT  19.100 155.140 19.420 171.290 ;
        RECT  53.655 155.035 53.935 171.290 ;
        RECT  56.365 155.280 56.645 171.315 ;
        RECT  57.120 155.300 57.400 171.315 ;
        RECT  57.835 155.130 58.115 171.315 ;
        RECT  0.600 155.310 64.400 171.290 ;
        RECT  56.240 155.310 61.880 171.315 ;
        RECT  53.895 155.310 55.870 171.370 ;
        RECT  31.880 155.310 32.380 171.375 ;
        RECT  3.210 155.310 3.490 171.380 ;
        RECT  34.655 155.310 38.715 171.480 ;
        RECT  39.605 155.310 42.020 171.480 ;
        RECT  2.000 0.000 63.000 60.210 ;
        RECT  0.600 0.600 64.400 60.210 ;
        RECT  0.600 0.600 1.210 135.520 ;
        RECT  0.600 91.020 64.400 135.520 ;
        RECT  4.080 91.020 60.940 135.690 ;
        RECT  62.580 91.020 62.995 135.710 ;
        LAYER M3 ;
        RECT  0.600 247.660 23.220 248.740 ;
        RECT  0.600 247.660 22.900 249.400 ;
        RECT  26.260 247.660 64.400 248.740 ;
        RECT  26.580 247.660 27.000 249.400 ;
        RECT  31.470 247.660 64.400 249.400 ;
        RECT  0.600 124.090 64.400 129.850 ;
        RECT  3.990 123.970 60.900 135.790 ;
        RECT  1.640 124.090 63.600 135.790 ;
        RECT  1.810 124.090 2.830 154.520 ;
        RECT  5.155 123.970 60.900 171.560 ;
        RECT  1.640 155.040 63.600 171.560 ;
        RECT  1.640 183.580 63.600 185.950 ;
        RECT  5.490 124.090 63.600 200.820 ;
        RECT  1.640 196.170 63.600 200.820 ;
        RECT  56.300 123.970 56.580 201.060 ;
        RECT  0.600 0.600 64.400 60.480 ;
        RECT  2.000 0.000 63.000 88.700 ;
        RECT  0.600 0.600 1.480 91.220 ;
        RECT  0.600 90.750 64.400 91.220 ;
        LAYER TOP_M ;
        RECT  0.600 247.690 64.400 248.850 ;
        RECT  0.600 247.690 23.010 249.400 ;
        RECT  26.470 247.690 27.110 249.400 ;
        RECT  31.360 247.690 64.400 249.400 ;
        RECT  2.000 0.000 63.000 91.190 ;
        RECT  0.600 0.600 64.400 91.190 ;
    END
END pc3b01u

MACRO pc3b01d
    CLASS PAD ;
    FOREIGN pc3b01d 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 65.000 BY 250.000 ;
    SYMMETRY X Y R90 ;
    SITE IOSite_c ;
    PIN PAD
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 55.440  LAYER TOP_M  ;
        ANTENNAPARTIALMETALSIDEAREA 287.938  LAYER M3  ;
        ANTENNAPARTIALMETALSIDEAREA 480.740  LAYER M2  ;
        ANTENNADIFFAREA 2657.280  LAYER TOP_M  ;
        ANTENNADIFFAREA 2657.280  LAYER M3  ;
        ANTENNADIFFAREA 1209.600  LAYER M2  ;
        ANTENNAPARTIALCUTAREA 632.318  LAYER TOP_V  ;
        ANTENNAPARTIALCUTAREA 349.898  LAYER V3  ;
        ANTENNAPARTIALCUTAREA 255.798  LAYER V2  ;
        PORT
        LAYER M3 ;
        RECT  23.740 249.580 25.740 250.000 ;
        LAYER M2 ;
        RECT  2.000 61.000 63.000 90.230 ;
        RECT  23.740 246.275 25.740 250.000 ;
        END
    END PAD
    PIN OEN
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 67.374  LAYER M1  ;
        ANTENNAPARTIALMETALSIDEAREA 80.634  LAYER M2  ;
        ANTENNAPARTIALMETALSIDEAREA 41.679  LAYER M3  ;
        ANTENNADIFFAREA 0.250  LAYER M3  ;
        ANTENNAPARTIALCUTAREA 0.203  LAYER V2  ;
        ANTENNAPARTIALCUTAREA 0.135  LAYER V3  ;
        ANTENNAGATEAREA 8.100  LAYER M2  ;
        ANTENNAGATEAREA 9.900  LAYER M3  ;
        PORT
        LAYER M3 ;
        RECT  29.900 249.580 30.630 250.000 ;
        LAYER M2 ;
        RECT  29.900 249.580 30.630 250.000 ;
        END
    END OEN
    PIN CIN
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 32.277  LAYER M3  ;
        ANTENNAPARTIALMETALSIDEAREA 96.916  LAYER M2  ;
        ANTENNAPARTIALMETALSIDEAREA 67.374  LAYER M1  ;
        ANTENNADIFFAREA 20.600  LAYER M3  ;
        ANTENNAPARTIALCUTAREA 0.135  LAYER V3  ;
        ANTENNAPARTIALCUTAREA 0.203  LAYER V2  ;
        PORT
        LAYER M3 ;
        RECT  28.870 249.580 29.600 250.000 ;
        LAYER M2 ;
        RECT  28.870 249.580 29.600 250.000 ;
        END
    END CIN
    PIN I
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 80.804  LAYER M2  ;
        ANTENNAPARTIALMETALSIDEAREA 67.374  LAYER M1  ;
        ANTENNAPARTIALMETALSIDEAREA 41.096  LAYER M3  ;
        ANTENNADIFFAREA 0.250  LAYER M3  ;
        ANTENNAPARTIALCUTAREA 0.203  LAYER V2  ;
        ANTENNAPARTIALCUTAREA 0.135  LAYER V3  ;
        ANTENNAGATEAREA 8.100  LAYER M2  ;
        ANTENNAGATEAREA 9.900  LAYER M3  ;
        PORT
        LAYER M3 ;
        RECT  27.840 249.580 28.570 250.000 ;
        LAYER M2 ;
        RECT  27.840 249.580 28.570 250.000 ;
        END
    END I
    PIN VDDO
        DIRECTION INOUT ;
        USE power ;
        PORT
        LAYER M3 ;
        RECT  64.200 192.330 65.000 200.640 ;
        RECT  0.000 201.660 65.000 221.520 ;
        RECT  0.000 222.720 65.000 246.820 ;
        RECT  0.000 192.330 0.800 200.640 ;
        LAYER M2 ;
        RECT  0.000 186.470 65.000 195.650 ;
        LAYER TOP_M ;
        RECT  0.000 195.170 65.000 200.640 ;
        RECT  0.000 201.660 65.000 221.520 ;
        RECT  0.000 222.720 65.000 246.820 ;
        END
    END VDDO
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        PORT
        LAYER M3 ;
        RECT  64.200 163.510 65.000 190.890 ;
        RECT  0.000 163.510 0.800 190.890 ;
        LAYER M2 ;
        RECT  0.000 172.080 65.000 183.060 ;
        LAYER TOP_M ;
        RECT  0.000 163.500 65.000 194.560 ;
        END
    END VDD
    PIN VSSO
        DIRECTION INOUT ;
        USE ground ;
        PORT
        LAYER M3 ;
        RECT  0.000 92.060 65.000 123.250 ;
        RECT  64.200 149.940 65.000 162.610 ;
        RECT  0.000 149.940 0.800 162.610 ;
        LAYER M2 ;
        RECT  0.000 147.040 65.000 154.520 ;
        LAYER TOP_M ;
        RECT  0.000 92.060 65.000 123.250 ;
        RECT  0.000 155.410 65.000 162.610 ;
        END
    END VSSO
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        PORT
        LAYER M3 ;
        RECT  64.200 130.690 65.000 148.880 ;
        RECT  0.000 130.690 0.800 148.880 ;
        LAYER M2 ;
        RECT  0.000 136.310 65.000 146.340 ;
        LAYER TOP_M ;
        RECT  0.000 123.850 65.000 154.560 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  2.000 0.000 63.000 250.000 ;
        RECT  0.000 88.990 65.000 130.360 ;
        RECT  0.000 136.510 65.000 157.550 ;
        RECT  0.315 158.150 64.700 158.460 ;
        RECT  0.300 158.930 64.700 159.230 ;
        RECT  0.300 159.530 64.700 159.830 ;
        RECT  0.300 160.130 64.700 160.430 ;
        RECT  0.300 160.730 64.700 161.030 ;
        RECT  0.300 161.330 64.700 161.630 ;
        RECT  0.300 161.910 64.700 162.190 ;
        RECT  0.300 162.490 64.700 162.770 ;
        RECT  0.300 163.070 64.700 163.350 ;
        RECT  0.300 163.650 64.700 163.950 ;
        RECT  0.300 164.250 64.700 164.550 ;
        RECT  0.300 164.850 64.700 165.150 ;
        RECT  0.300 165.450 64.700 165.750 ;
        RECT  0.300 166.050 64.700 166.350 ;
        RECT  0.300 166.650 64.700 166.960 ;
        RECT  0.300 167.260 64.700 167.560 ;
        RECT  0.300 167.860 64.700 168.160 ;
        RECT  0.000 169.150 65.000 197.240 ;
        RECT  0.600 0.600 64.400 250.000 ;
        RECT  0.000 198.470 65.000 250.000 ;
        LAYER M2 ;
        RECT  1.840 196.420 2.120 249.400 ;
        RECT  63.180 196.430 63.670 249.400 ;
        RECT  0.600 196.440 64.400 245.485 ;
        RECT  26.530 196.440 64.400 248.790 ;
        RECT  0.600 196.440 22.950 249.400 ;
        RECT  26.530 196.440 27.050 249.400 ;
        RECT  31.420 196.440 64.400 249.400 ;
        RECT  14.290 183.720 52.380 185.680 ;
        RECT  0.600 183.850 64.400 185.680 ;
        RECT  54.910 183.850 57.160 185.865 ;
        RECT  46.230 183.720 51.730 185.870 ;
        RECT  18.450 155.160 18.800 171.290 ;
        RECT  19.100 155.140 19.420 171.290 ;
        RECT  49.250 155.125 51.490 171.290 ;
        RECT  52.430 155.295 52.740 171.290 ;
        RECT  53.655 155.035 53.935 171.290 ;
        RECT  56.365 155.280 56.645 171.315 ;
        RECT  57.120 155.300 57.400 171.315 ;
        RECT  57.835 155.130 58.115 171.315 ;
        RECT  0.600 155.310 64.400 171.290 ;
        RECT  56.240 155.310 61.880 171.315 ;
        RECT  53.895 155.310 55.870 171.370 ;
        RECT  3.210 155.310 3.490 171.380 ;
        RECT  34.655 155.310 38.715 171.480 ;
        RECT  39.605 155.310 42.020 171.480 ;
        RECT  2.000 0.000 63.000 60.210 ;
        RECT  0.600 0.600 64.400 60.210 ;
        RECT  0.600 0.600 1.210 135.520 ;
        RECT  0.600 91.020 64.400 135.520 ;
        RECT  4.080 91.020 60.940 135.690 ;
        RECT  62.580 91.020 62.995 135.710 ;
        LAYER M3 ;
        RECT  0.600 247.660 23.220 248.740 ;
        RECT  0.600 247.660 22.900 249.400 ;
        RECT  26.260 247.660 64.400 248.740 ;
        RECT  26.580 247.660 27.000 249.400 ;
        RECT  31.470 247.660 64.400 249.400 ;
        RECT  0.600 124.090 64.400 129.850 ;
        RECT  3.990 123.970 60.900 135.790 ;
        RECT  1.640 124.090 63.600 135.790 ;
        RECT  1.810 124.090 2.830 154.520 ;
        RECT  5.155 123.970 60.900 171.560 ;
        RECT  1.640 155.040 63.600 171.560 ;
        RECT  1.640 183.580 63.600 185.950 ;
        RECT  5.490 124.090 63.600 200.820 ;
        RECT  1.640 196.170 63.600 200.820 ;
        RECT  56.300 123.970 56.580 201.060 ;
        RECT  0.600 0.600 64.400 60.480 ;
        RECT  2.000 0.000 63.000 88.700 ;
        RECT  0.600 0.600 1.480 91.220 ;
        RECT  0.600 90.750 64.400 91.220 ;
        LAYER TOP_M ;
        RECT  0.600 247.690 64.400 248.850 ;
        RECT  0.600 247.690 23.010 249.400 ;
        RECT  26.470 247.690 27.110 249.400 ;
        RECT  31.360 247.690 64.400 249.400 ;
        RECT  2.000 0.000 63.000 91.190 ;
        RECT  0.600 0.600 64.400 91.190 ;
    END
END pc3b01d

MACRO pc3b01
    CLASS PAD ;
    FOREIGN pc3b01 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 65.000 BY 250.000 ;
    SYMMETRY X Y R90 ;
    SITE IOSite_c ;
    PIN PAD
        DIRECTION INOUT ;
        ANTENNAPARTIALMETALSIDEAREA 55.440  LAYER TOP_M  ;
        ANTENNAPARTIALMETALSIDEAREA 287.938  LAYER M3  ;
        ANTENNAPARTIALMETALSIDEAREA 480.740  LAYER M2  ;
        ANTENNADIFFAREA 2657.280  LAYER TOP_M  ;
        ANTENNADIFFAREA 2657.280  LAYER M3  ;
        ANTENNADIFFAREA 1209.600  LAYER M2  ;
        ANTENNAPARTIALCUTAREA 632.318  LAYER TOP_V  ;
        ANTENNAPARTIALCUTAREA 349.898  LAYER V3  ;
        ANTENNAPARTIALCUTAREA 255.798  LAYER V2  ;
        PORT
        LAYER M3 ;
        RECT  23.740 249.580 25.740 250.000 ;
        LAYER M2 ;
        RECT  2.000 61.000 63.000 90.230 ;
        RECT  23.740 246.275 25.740 250.000 ;
        END
    END PAD
    PIN OEN
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 67.374  LAYER M1  ;
        ANTENNAPARTIALMETALSIDEAREA 80.634  LAYER M2  ;
        ANTENNAPARTIALMETALSIDEAREA 41.679  LAYER M3  ;
        ANTENNADIFFAREA 0.250  LAYER M3  ;
        ANTENNAPARTIALCUTAREA 0.203  LAYER V2  ;
        ANTENNAPARTIALCUTAREA 0.135  LAYER V3  ;
        ANTENNAGATEAREA 8.100  LAYER M2  ;
        ANTENNAGATEAREA 9.900  LAYER M3  ;
        PORT
        LAYER M3 ;
        RECT  29.900 249.580 30.630 250.000 ;
        LAYER M2 ;
        RECT  29.900 249.580 30.630 250.000 ;
        END
    END OEN
    PIN CIN
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 32.277  LAYER M3  ;
        ANTENNAPARTIALMETALSIDEAREA 96.916  LAYER M2  ;
        ANTENNAPARTIALMETALSIDEAREA 67.374  LAYER M1  ;
        ANTENNADIFFAREA 20.600  LAYER M3  ;
        ANTENNAPARTIALCUTAREA 0.135  LAYER V3  ;
        ANTENNAPARTIALCUTAREA 0.203  LAYER V2  ;
        PORT
        LAYER M3 ;
        RECT  28.870 249.580 29.600 250.000 ;
        LAYER M2 ;
        RECT  28.870 249.580 29.600 250.000 ;
        END
    END CIN
    PIN I
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 80.804  LAYER M2  ;
        ANTENNAPARTIALMETALSIDEAREA 67.374  LAYER M1  ;
        ANTENNAPARTIALMETALSIDEAREA 41.096  LAYER M3  ;
        ANTENNADIFFAREA 0.250  LAYER M3  ;
        ANTENNAPARTIALCUTAREA 0.203  LAYER V2  ;
        ANTENNAPARTIALCUTAREA 0.135  LAYER V3  ;
        ANTENNAGATEAREA 8.100  LAYER M2  ;
        ANTENNAGATEAREA 9.900  LAYER M3  ;
        PORT
        LAYER M3 ;
        RECT  27.840 249.580 28.570 250.000 ;
        LAYER M2 ;
        RECT  27.840 249.580 28.570 250.000 ;
        END
    END I
    PIN VDDO
        DIRECTION INOUT ;
        USE power ;
        PORT
        LAYER M3 ;
        RECT  64.200 192.330 65.000 200.640 ;
        RECT  0.000 201.660 65.000 221.520 ;
        RECT  0.000 222.720 65.000 246.820 ;
        RECT  0.000 192.330 0.800 200.640 ;
        LAYER M2 ;
        RECT  0.000 186.470 65.000 195.650 ;
        LAYER TOP_M ;
        RECT  0.000 195.170 65.000 200.640 ;
        RECT  0.000 201.660 65.000 221.520 ;
        RECT  0.000 222.720 65.000 246.820 ;
        END
    END VDDO
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        PORT
        LAYER M3 ;
        RECT  64.200 163.510 65.000 190.890 ;
        RECT  0.000 163.510 0.800 190.890 ;
        LAYER M2 ;
        RECT  0.000 172.080 65.000 183.060 ;
        LAYER TOP_M ;
        RECT  0.000 163.500 65.000 194.560 ;
        END
    END VDD
    PIN VSSO
        DIRECTION INOUT ;
        USE ground ;
        PORT
        LAYER M3 ;
        RECT  0.000 92.060 65.000 123.250 ;
        RECT  64.200 149.940 65.000 162.610 ;
        RECT  0.000 149.940 0.800 162.610 ;
        LAYER M2 ;
        RECT  0.000 147.040 65.000 154.520 ;
        LAYER TOP_M ;
        RECT  0.000 92.060 65.000 123.250 ;
        RECT  0.000 155.410 65.000 162.610 ;
        END
    END VSSO
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        PORT
        LAYER M3 ;
        RECT  64.200 130.690 65.000 148.880 ;
        RECT  0.000 130.690 0.800 148.880 ;
        LAYER M2 ;
        RECT  0.000 136.310 65.000 146.340 ;
        LAYER TOP_M ;
        RECT  0.000 123.850 65.000 154.560 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  2.000 0.000 63.000 250.000 ;
        RECT  0.000 88.990 65.000 130.360 ;
        RECT  0.000 136.510 65.000 157.550 ;
        RECT  0.315 158.150 64.700 158.460 ;
        RECT  0.300 158.930 64.700 159.230 ;
        RECT  0.300 159.530 64.700 159.830 ;
        RECT  0.300 160.130 64.700 160.430 ;
        RECT  0.300 160.730 64.700 161.030 ;
        RECT  0.300 161.330 64.700 161.630 ;
        RECT  0.300 161.910 64.700 162.190 ;
        RECT  0.300 162.490 64.700 162.770 ;
        RECT  0.300 163.070 64.700 163.350 ;
        RECT  0.300 163.650 64.700 163.950 ;
        RECT  0.300 164.250 64.700 164.550 ;
        RECT  0.300 164.850 64.700 165.150 ;
        RECT  0.300 165.450 64.700 165.750 ;
        RECT  0.300 166.050 64.700 166.350 ;
        RECT  0.300 166.650 64.700 166.960 ;
        RECT  0.300 167.260 64.700 167.560 ;
        RECT  0.300 167.860 64.700 168.160 ;
        RECT  0.000 169.150 65.000 197.240 ;
        RECT  0.600 0.600 64.400 250.000 ;
        RECT  0.000 198.470 65.000 250.000 ;
        LAYER M2 ;
        RECT  1.840 196.420 2.120 249.400 ;
        RECT  63.180 196.430 63.670 249.400 ;
        RECT  0.600 196.440 64.400 245.485 ;
        RECT  26.530 196.440 64.400 248.790 ;
        RECT  0.600 196.440 22.950 249.400 ;
        RECT  26.530 196.440 27.050 249.400 ;
        RECT  31.420 196.440 64.400 249.400 ;
        RECT  14.290 183.720 52.380 185.680 ;
        RECT  0.600 183.850 64.400 185.680 ;
        RECT  54.910 183.850 57.160 185.865 ;
        RECT  46.230 183.720 51.730 185.870 ;
        RECT  18.450 155.160 18.800 171.290 ;
        RECT  19.100 155.140 19.420 171.290 ;
        RECT  53.655 155.035 53.935 171.290 ;
        RECT  56.365 155.280 56.645 171.315 ;
        RECT  57.120 155.300 57.400 171.315 ;
        RECT  57.835 155.130 58.115 171.315 ;
        RECT  0.600 155.310 64.400 171.290 ;
        RECT  56.240 155.310 61.880 171.315 ;
        RECT  53.895 155.310 55.870 171.370 ;
        RECT  3.210 155.310 3.490 171.380 ;
        RECT  34.655 155.310 38.715 171.480 ;
        RECT  39.605 155.310 42.020 171.480 ;
        RECT  2.000 0.000 63.000 60.210 ;
        RECT  0.600 0.600 64.400 60.210 ;
        RECT  0.600 0.600 1.210 135.520 ;
        RECT  0.600 91.020 64.400 135.520 ;
        RECT  4.080 91.020 60.940 135.690 ;
        RECT  62.580 91.020 62.995 135.710 ;
        LAYER M3 ;
        RECT  0.600 247.660 23.220 248.740 ;
        RECT  0.600 247.660 22.900 249.400 ;
        RECT  26.260 247.660 64.400 248.740 ;
        RECT  26.580 247.660 27.000 249.400 ;
        RECT  31.470 247.660 64.400 249.400 ;
        RECT  0.600 124.090 64.400 129.850 ;
        RECT  3.990 123.970 60.900 135.790 ;
        RECT  1.640 124.090 63.600 135.790 ;
        RECT  1.810 124.090 2.830 154.520 ;
        RECT  5.155 123.970 60.900 171.560 ;
        RECT  1.640 155.040 63.600 171.560 ;
        RECT  1.640 183.580 63.600 185.950 ;
        RECT  5.490 124.090 63.600 200.820 ;
        RECT  1.640 196.170 63.600 200.820 ;
        RECT  56.300 123.970 56.580 201.060 ;
        RECT  0.600 0.600 64.400 60.480 ;
        RECT  2.000 0.000 63.000 88.700 ;
        RECT  0.600 0.600 1.480 91.220 ;
        RECT  0.600 90.750 64.400 91.220 ;
        LAYER TOP_M ;
        RECT  0.600 247.690 64.400 248.850 ;
        RECT  0.600 247.690 23.010 249.400 ;
        RECT  26.470 247.690 27.110 249.400 ;
        RECT  31.360 247.690 64.400 249.400 ;
        RECT  2.000 0.000 63.000 91.190 ;
        RECT  0.600 0.600 64.400 91.190 ;
    END
END pc3b01

MACRO apvdi
    CLASS PAD ;
    FOREIGN apvdi 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 65.000 BY 250.000 ;
    SYMMETRY X Y R90 ;
    SITE IOSite_c ;
    PIN AVSSO
        DIRECTION INOUT ;
        USE ground ;
        PORT
        LAYER M3 ;
        RECT  0.000 92.060 65.000 123.250 ;
        RECT  64.200 149.940 65.000 162.610 ;
        RECT  0.000 149.940 0.800 162.610 ;
        LAYER M2 ;
        RECT  0.000 147.040 65.000 154.520 ;
        LAYER TOP_M ;
        RECT  0.000 92.060 65.000 123.250 ;
        RECT  0.000 155.410 65.000 162.610 ;
        END
    END AVSSO
    PIN AVSS
        DIRECTION INOUT ;
        USE ground ;
        PORT
        LAYER M3 ;
        RECT  64.200 141.450 65.000 148.880 ;
        RECT  0.000 141.450 0.800 148.880 ;
        LAYER M2 ;
        RECT  0.000 143.070 65.000 146.340 ;
        RECT  57.840 136.310 65.000 146.340 ;
        RECT  0.000 136.310 6.265 146.340 ;
        LAYER TOP_M ;
        RECT  0.000 141.450 65.000 154.560 ;
        END
    END AVSS
    PIN AVDD
        DIRECTION OUTPUT ;
        USE power ;
        PORT
	CLASS CORE ;
        LAYER M3 ;
        RECT  64.200 163.510 65.000 190.890 ;
        RECT  15.560 247.440 49.380 250.000 ;
        RECT  0.000 163.510 0.800 190.890 ;
        LAYER M2 ;
        RECT  0.000 172.080 65.000 183.060 ;
        RECT  2.000 61.000 63.000 90.230 ;
        RECT  15.560 242.060 49.380 250.000 ;
        LAYER TOP_M ;
        RECT  0.000 163.500 65.000 194.560 ;
        RECT  15.560 247.440 49.380 250.000 ;
        END
    END AVDD
    PIN AVDDO
        DIRECTION INOUT ;
        USE power ;
        PORT
        LAYER M3 ;
        RECT  64.200 192.330 65.000 200.640 ;
        RECT  0.000 201.660 65.000 218.520 ;
        RECT  0.000 219.720 65.000 246.820 ;
        RECT  0.000 192.330 0.800 200.640 ;
        LAYER M2 ;
        RECT  0.000 186.470 65.000 194.870 ;
        LAYER TOP_M ;
        RECT  0.000 195.170 65.000 200.640 ;
        RECT  0.000 201.660 65.000 221.520 ;
        RECT  0.000 222.720 65.000 246.820 ;
        END
    END AVDDO
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        PORT
        LAYER M3 ;
        RECT  64.200 130.680 65.000 140.840 ;
        RECT  0.000 130.680 0.800 140.840 ;
        LAYER TOP_M ;
        RECT  0.000 123.850 65.000 140.850 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  2.000 0.000 63.000 249.570 ;
        RECT  0.000 88.990 65.000 130.360 ;
        RECT  0.000 136.510 65.000 157.550 ;
        RECT  0.500 136.510 64.500 160.550 ;
        RECT  0.000 192.990 65.000 194.230 ;
        RECT  0.000 195.470 65.000 247.000 ;
        RECT  0.600 0.600 64.400 249.570 ;
        RECT  0.000 248.330 65.000 249.570 ;
        LAYER M2 ;
        RECT  50.010 195.470 52.110 241.270 ;
        RECT  0.600 195.660 64.400 241.270 ;
        RECT  12.630 195.470 14.950 243.720 ;
        RECT  50.060 195.660 64.400 243.720 ;
        RECT  0.600 195.660 14.770 249.400 ;
        RECT  50.170 195.660 64.400 249.400 ;
        RECT  0.780 195.660 6.550 249.570 ;
        RECT  0.600 183.850 64.400 185.680 ;
        RECT  0.600 155.310 64.400 171.290 ;
        RECT  2.000 0.000 63.000 60.210 ;
        RECT  0.600 0.600 64.400 60.210 ;
        RECT  0.600 0.600 1.210 135.520 ;
        RECT  0.600 91.020 64.400 135.520 ;
        RECT  4.080 91.020 60.940 135.690 ;
        RECT  7.055 91.020 57.050 142.470 ;
        RECT  7.025 136.310 57.155 142.470 ;
        LAYER M3 ;
        RECT  0.600 247.660 14.720 249.400 ;
        RECT  0.775 247.660 6.560 249.570 ;
        RECT  50.220 247.660 64.400 249.400 ;
        RECT  0.600 124.090 64.400 129.840 ;
        RECT  1.400 124.090 63.360 135.790 ;
        RECT  62.175 124.090 63.250 154.300 ;
        RECT  1.400 124.090 2.850 154.470 ;
        RECT  3.530 124.090 59.560 200.820 ;
        RECT  60.380 136.230 61.520 200.820 ;
        RECT  1.640 155.040 63.360 171.560 ;
        RECT  1.640 183.580 63.360 185.950 ;
        RECT  3.530 155.040 63.255 200.820 ;
        RECT  1.640 195.390 63.360 200.820 ;
        RECT  62.175 155.040 63.255 200.960 ;
        RECT  58.475 155.040 60.775 201.060 ;
        RECT  0.600 0.600 64.400 60.480 ;
        RECT  2.000 0.000 63.000 88.700 ;
        RECT  0.600 0.600 1.480 91.220 ;
        RECT  0.600 90.750 64.400 91.220 ;
        LAYER TOP_M ;
        RECT  0.600 247.690 14.690 249.400 ;
        RECT  50.250 247.690 64.400 249.400 ;
        RECT  2.000 0.000 63.000 91.190 ;
        RECT  0.600 0.600 64.400 91.190 ;
    END
END apvdi

MACRO apvda
    CLASS PAD ;
    FOREIGN apvda 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 65.000 BY 250.000 ;
    SYMMETRY X Y R90 ;
    SITE IOSite_c ;
    PIN AVSSO
        DIRECTION INOUT ;
        USE ground ;
        PORT
        LAYER M3 ;
        RECT  64.200 92.060 65.000 123.250 ;
        RECT  0.000 92.060 65.000 122.850 ;
        RECT  0.000 92.060 2.850 123.250 ;
        RECT  64.200 149.940 65.000 162.610 ;
        RECT  0.000 149.940 0.800 162.610 ;
        LAYER M2 ;
        RECT  0.000 147.040 65.000 154.520 ;
        LAYER TOP_M ;
        RECT  0.000 92.060 65.000 123.250 ;
        RECT  0.000 155.410 65.000 162.610 ;
        END
    END AVSSO
    PIN AVSS
        DIRECTION INOUT ;
        USE ground ;
        PORT
        LAYER M3 ;
        RECT  64.200 141.450 65.000 148.880 ;
        RECT  0.000 141.450 0.800 148.880 ;
        LAYER M2 ;
        RECT  0.000 143.070 65.000 146.340 ;
        RECT  57.840 136.310 65.000 146.340 ;
        RECT  0.000 136.310 6.265 146.340 ;
        LAYER TOP_M ;
        RECT  0.000 141.450 65.000 154.560 ;
        END
    END AVSS
    PIN AVDD
        DIRECTION INOUT ;
        USE power ;
        PORT
        LAYER M3 ;
        RECT  64.200 163.510 65.000 190.890 ;
        RECT  0.000 163.510 0.800 190.890 ;
        LAYER M2 ;
        RECT  0.000 172.080 65.000 183.060 ;
        LAYER TOP_M ;
        RECT  0.000 163.500 65.000 194.560 ;
        END
    END AVDD
    PIN AVDDO
        DIRECTION OUTPUT ;
        USE power ;
        PORT
        LAYER M3 ;
        RECT  64.200 192.330 65.000 200.640 ;
        RECT  0.000 201.660 65.000 218.520 ;
        RECT  0.000 219.720 65.000 246.820 ;
        RECT  0.000 192.330 0.800 200.640 ;
        LAYER M2 ;
        RECT  0.000 186.470 65.000 194.870 ;
        RECT  2.000 61.000 63.000 90.230 ;
        LAYER TOP_M ;
        RECT  0.000 195.170 65.000 200.640 ;
        RECT  0.000 201.660 65.000 221.520 ;
        RECT  0.000 222.720 65.000 246.820 ;
        END
    END AVDDO
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        PORT
        LAYER M3 ;
        RECT  64.200 130.680 65.000 140.840 ;
        RECT  0.000 130.680 0.800 140.840 ;
        LAYER TOP_M ;
        RECT  0.000 123.850 65.000 140.850 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  2.000 0.000 63.000 249.570 ;
        RECT  0.000 88.990 65.000 130.360 ;
        RECT  0.000 136.510 65.000 157.550 ;
        RECT  0.500 136.510 64.500 160.550 ;
        RECT  0.000 192.990 65.000 194.230 ;
        RECT  0.000 195.470 65.000 247.000 ;
        RECT  0.600 0.600 64.400 249.570 ;
        RECT  0.000 248.330 65.000 249.570 ;
        LAYER M2 ;
        RECT  12.640 195.470 14.730 249.400 ;
        RECT  50.010 195.470 52.020 249.400 ;
        RECT  0.600 195.660 64.400 249.400 ;
        RECT  0.780 195.660 6.550 249.570 ;
        RECT  0.600 183.850 64.400 185.680 ;
        RECT  0.600 155.310 64.400 171.290 ;
        RECT  2.000 0.000 63.000 60.210 ;
        RECT  0.600 0.600 64.400 60.210 ;
        RECT  0.600 0.600 1.210 135.520 ;
        RECT  0.600 91.020 64.400 135.520 ;
        RECT  4.080 91.020 60.940 135.690 ;
        RECT  7.055 91.020 57.050 142.470 ;
        RECT  7.025 136.310 57.155 142.470 ;
        LAYER M3 ;
        RECT  0.600 247.660 64.400 249.400 ;
        RECT  0.775 247.660 6.560 249.570 ;
        RECT  0.600 124.090 64.400 129.840 ;
        RECT  3.690 123.690 63.360 135.790 ;
        RECT  1.400 124.090 63.360 135.790 ;
        RECT  1.400 124.090 2.850 154.470 ;
        RECT  3.745 123.690 59.560 200.820 ;
        RECT  60.380 149.370 61.520 200.820 ;
        RECT  1.640 155.040 63.360 171.560 ;
        RECT  1.640 183.580 63.360 185.950 ;
        RECT  3.745 155.040 63.255 200.820 ;
        RECT  1.640 195.390 63.360 200.820 ;
        RECT  62.175 155.040 63.255 200.960 ;
        RECT  7.270 123.690 9.370 201.060 ;
        RECT  55.630 123.690 57.730 201.060 ;
        RECT  58.475 155.040 60.775 201.060 ;
        RECT  0.600 0.600 64.400 60.480 ;
        RECT  2.000 0.000 63.000 88.700 ;
        RECT  0.600 0.600 1.480 91.220 ;
        RECT  0.600 90.750 64.400 91.220 ;
        LAYER TOP_M ;
        RECT  0.600 247.690 64.400 249.400 ;
        RECT  2.000 0.000 63.000 91.190 ;
        RECT  0.600 0.600 64.400 91.190 ;
    END
END apvda

MACRO apv0i
    CLASS PAD ;
    FOREIGN apv0i 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 65.000 BY 250.000 ;
    SYMMETRY X Y R90 ;
    SITE IOSite_c ;
    PIN AVSSO
        DIRECTION INOUT ;
        USE ground ;
        PORT
        LAYER M3 ;
        RECT  62.810 92.060 65.000 123.250 ;
        RECT  0.000 92.060 65.000 118.650 ;
        RECT  0.000 92.060 2.850 123.250 ;
        RECT  64.200 149.940 65.000 162.610 ;
        RECT  0.000 149.940 0.800 162.610 ;
        LAYER M2 ;
        RECT  0.000 147.040 65.000 154.520 ;
        LAYER TOP_M ;
        RECT  0.000 92.060 65.000 123.250 ;
        RECT  0.000 155.410 65.000 162.610 ;
        END
    END AVSSO
    PIN AVSS
        DIRECTION OUTPUT ;
        USE ground ;
        PORT
	CLASS CORE ;
        LAYER M3 ;
        RECT  64.200 141.450 65.000 148.880 ;
        RECT  15.570 247.420 49.400 250.000 ;
        RECT  0.000 141.450 0.800 148.880 ;
        LAYER M2 ;
        RECT  0.000 143.070 65.000 146.340 ;
        RECT  57.840 136.310 65.000 146.340 ;
        RECT  0.000 136.310 6.265 146.340 ;
        RECT  2.000 61.000 63.000 90.230 ;
        RECT  15.560 243.630 49.380 250.000 ;
        LAYER TOP_M ;
        RECT  0.000 141.450 65.000 154.560 ;
        RECT  15.560 247.420 49.380 250.000 ;
        END
    END AVSS
    PIN AVDD
        DIRECTION INOUT ;
        USE power ;
        PORT
        LAYER M3 ;
        RECT  64.200 163.510 65.000 190.890 ;
        RECT  0.000 163.510 0.800 190.890 ;
        LAYER M2 ;
        RECT  0.000 172.080 65.000 183.060 ;
        LAYER TOP_M ;
        RECT  0.000 163.500 65.000 194.560 ;
        END
    END AVDD
    PIN AVDDO
        DIRECTION INOUT ;
        USE power ;
        PORT
        LAYER M3 ;
        RECT  64.200 192.330 65.000 200.640 ;
        RECT  0.000 201.660 65.000 218.520 ;
        RECT  0.000 219.720 65.000 246.820 ;
        RECT  0.000 192.330 0.800 200.640 ;
        LAYER M2 ;
        RECT  0.000 186.470 65.000 194.870 ;
        LAYER TOP_M ;
        RECT  0.000 195.170 65.000 200.640 ;
        RECT  0.000 201.660 65.000 221.520 ;
        RECT  0.000 222.720 65.000 246.820 ;
        END
    END AVDDO
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        PORT
        LAYER M3 ;
        RECT  64.200 130.680 65.000 140.840 ;
        RECT  0.000 130.680 0.800 140.840 ;
        LAYER TOP_M ;
        RECT  0.000 123.850 65.000 140.850 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  2.000 0.000 63.000 249.570 ;
        RECT  0.000 88.990 65.000 130.360 ;
        RECT  0.000 136.510 65.000 157.550 ;
        RECT  0.500 136.510 64.500 160.550 ;
        RECT  0.000 192.990 65.000 194.230 ;
        RECT  0.000 195.470 65.000 247.000 ;
        RECT  0.600 0.600 64.400 249.570 ;
        RECT  0.000 248.330 65.000 249.570 ;
        LAYER M2 ;
        RECT  12.640 195.470 14.730 249.400 ;
        RECT  50.010 195.470 52.020 242.840 ;
        RECT  0.600 195.660 64.400 242.840 ;
        RECT  0.600 195.660 14.950 243.720 ;
        RECT  50.060 195.660 64.400 243.720 ;
        RECT  0.600 195.660 14.770 249.400 ;
        RECT  50.170 195.660 64.400 249.400 ;
        RECT  0.780 195.660 6.550 249.570 ;
        RECT  0.600 183.850 64.400 185.680 ;
        RECT  0.600 155.310 64.400 171.290 ;
        RECT  2.000 0.000 63.000 60.210 ;
        RECT  0.600 0.600 64.400 60.210 ;
        RECT  0.600 0.600 1.210 135.520 ;
        RECT  0.600 91.020 64.400 135.520 ;
        RECT  1.760 91.020 63.020 135.690 ;
        RECT  7.055 91.020 57.050 142.470 ;
        RECT  7.025 136.310 57.155 142.470 ;
        LAYER M3 ;
        RECT  0.600 247.660 14.730 249.400 ;
        RECT  0.775 247.660 6.560 249.570 ;
        RECT  50.240 247.660 64.400 249.400 ;
        RECT  3.450 119.490 61.970 135.790 ;
        RECT  0.600 124.090 64.400 129.840 ;
        RECT  1.400 124.090 63.360 135.790 ;
        RECT  1.400 124.090 2.850 154.470 ;
        RECT  3.450 119.310 61.920 200.820 ;
        RECT  1.640 155.040 63.540 190.885 ;
        RECT  3.450 155.040 63.540 200.310 ;
        RECT  62.460 139.485 63.540 200.310 ;
        RECT  1.640 195.390 63.360 200.820 ;
        RECT  0.600 0.600 64.400 60.480 ;
        RECT  2.000 0.000 63.000 88.700 ;
        RECT  0.600 0.600 1.480 91.220 ;
        RECT  0.600 90.750 64.400 91.220 ;
        LAYER TOP_M ;
        RECT  0.600 247.690 14.690 249.400 ;
        RECT  50.250 247.690 64.400 249.400 ;
        RECT  2.000 0.000 63.000 91.190 ;
        RECT  0.600 0.600 64.400 91.190 ;
    END
END apv0i

MACRO apv0a
    CLASS PAD ;
    FOREIGN apv0a 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 65.000 BY 250.000 ;
    SYMMETRY X Y R90 ;
    SITE IOSite_c ;
    PIN AVSSO
        DIRECTION OUTPUT ;
        USE ground ;
        PORT
        LAYER M3 ;
        RECT  62.345 92.060 65.000 123.250 ;
        RECT  0.000 92.060 65.000 118.905 ;
        RECT  0.000 92.060 2.850 123.250 ;
        RECT  64.200 149.940 65.000 162.610 ;
        RECT  0.000 149.940 0.800 162.610 ;
        LAYER M2 ;
        RECT  0.000 147.040 65.000 154.520 ;
        RECT  2.000 61.000 63.000 90.230 ;
        LAYER TOP_M ;
        RECT  0.000 92.060 65.000 123.250 ;
        RECT  0.000 155.410 65.000 162.610 ;
        END
    END AVSSO
    PIN AVSS
        DIRECTION INOUT ;
        USE ground ;
        PORT
        LAYER M3 ;
        RECT  64.200 141.450 65.000 148.880 ;
        RECT  0.000 141.450 0.800 148.880 ;
        LAYER M2 ;
        RECT  0.000 143.070 65.000 146.340 ;
        RECT  57.840 136.310 65.000 146.340 ;
        RECT  0.000 136.310 6.265 146.340 ;
        LAYER TOP_M ;
        RECT  0.000 141.450 65.000 154.560 ;
        END
    END AVSS
    PIN AVDD
        DIRECTION INOUT ;
        USE power ;
        PORT
        LAYER M3 ;
        RECT  64.200 163.510 65.000 190.890 ;
        RECT  0.000 163.510 0.800 190.890 ;
        LAYER M2 ;
        RECT  0.000 172.080 65.000 183.060 ;
        LAYER TOP_M ;
        RECT  0.000 163.500 65.000 194.560 ;
        END
    END AVDD
    PIN AVDDO
        DIRECTION INOUT ;
        USE power ;
        PORT
        LAYER M3 ;
        RECT  64.200 192.330 65.000 200.640 ;
        RECT  0.000 201.660 65.000 218.520 ;
        RECT  0.000 219.720 65.000 246.820 ;
        RECT  0.000 192.330 0.800 200.640 ;
        LAYER M2 ;
        RECT  0.000 186.470 65.000 194.870 ;
        LAYER TOP_M ;
        RECT  0.000 195.170 65.000 200.640 ;
        RECT  0.000 201.660 65.000 221.520 ;
        RECT  0.000 222.720 65.000 246.820 ;
        END
    END AVDDO
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        PORT
        LAYER M3 ;
        RECT  64.200 130.680 65.000 140.840 ;
        RECT  0.000 130.680 0.800 140.840 ;
        LAYER TOP_M ;
        RECT  0.000 123.850 65.000 140.850 ;
        END
    END VSS
    OBS
        LAYER M1 ;
        RECT  2.000 0.000 63.000 249.570 ;
        RECT  0.000 88.990 65.000 130.360 ;
        RECT  0.000 136.510 65.000 157.550 ;
        RECT  0.500 136.510 64.500 160.550 ;
        RECT  0.000 192.990 65.000 194.230 ;
        RECT  0.000 195.470 65.000 247.000 ;
        RECT  0.600 0.600 64.400 249.570 ;
        RECT  0.000 248.330 65.000 249.570 ;
        LAYER M2 ;
        RECT  12.640 195.470 14.730 249.400 ;
        RECT  50.010 195.470 52.020 249.400 ;
        RECT  0.600 195.660 64.400 249.400 ;
        RECT  0.780 195.660 6.550 249.570 ;
        RECT  0.600 183.850 64.400 185.680 ;
        RECT  0.600 155.310 64.400 171.290 ;
        RECT  2.000 0.000 63.000 60.210 ;
        RECT  0.600 0.600 64.400 60.210 ;
        RECT  0.600 0.600 1.210 135.520 ;
        RECT  0.600 91.020 64.400 135.520 ;
        RECT  1.970 91.020 63.080 135.690 ;
        RECT  7.055 91.020 57.050 142.470 ;
        RECT  7.025 136.310 57.155 142.470 ;
        LAYER M3 ;
        RECT  0.600 247.660 64.400 249.400 ;
        RECT  0.775 247.660 6.560 249.570 ;
        RECT  3.690 119.745 61.650 135.790 ;
        RECT  0.600 124.090 64.400 129.840 ;
        RECT  1.400 124.090 63.360 135.790 ;
        RECT  1.400 124.090 2.850 149.100 ;
        RECT  1.640 124.090 2.850 154.470 ;
        RECT  4.200 119.605 61.650 200.820 ;
        RECT  1.640 155.040 63.540 171.560 ;
        RECT  1.640 183.580 63.540 185.950 ;
        RECT  4.200 155.040 63.540 200.310 ;
        RECT  62.460 149.410 63.540 200.310 ;
        RECT  1.640 195.390 63.360 200.820 ;
        RECT  0.600 0.600 64.400 60.480 ;
        RECT  2.000 0.000 63.000 88.700 ;
        RECT  0.600 0.600 1.480 91.220 ;
        RECT  0.600 90.750 64.400 91.220 ;
        LAYER TOP_M ;
        RECT  0.600 247.690 64.400 249.400 ;
        RECT  2.000 0.000 63.000 91.190 ;
        RECT  0.600 0.600 64.400 91.190 ;
    END
END apv0a

MACRO apc3d01
    CLASS PAD ;
    FOREIGN apc3d01 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 65.000 BY 250.000 ;
    SYMMETRY X Y R90 ;
    SITE IOSite_c ;
    PIN PAD
        DIRECTION INPUT ;
        ANTENNAPARTIALMETALSIDEAREA 55.440  LAYER TOP_M  ;
        ANTENNAPARTIALMETALSIDEAREA 196.826  LAYER M3  ;
        ANTENNAPARTIALMETALSIDEAREA 480.740  LAYER M2  ;
        ANTENNADIFFAREA 2657.280  LAYER TOP_M  ;
        ANTENNADIFFAREA 2657.280  LAYER M3  ;
        ANTENNADIFFAREA 1209.600  LAYER M2  ;
        ANTENNAPARTIALCUTAREA 632.318  LAYER TOP_V  ;
        ANTENNAPARTIALCUTAREA 349.222  LAYER V3  ;
        ANTENNAPARTIALCUTAREA 255.798  LAYER V2  ;
        PORT
        LAYER M2 ;
        RECT  2.000 61.000 63.000 90.230 ;
        RECT  32.350 242.720 34.370 250.000 ;
        LAYER M3 ;
        RECT  32.350 249.580 34.370 250.000 ;
        END
    END PAD
    PIN CIN
        DIRECTION OUTPUT ;
        ANTENNAPARTIALMETALSIDEAREA 169.478  LAYER M2  ;
        ANTENNAPARTIALMETALSIDEAREA 67.374  LAYER M1  ;
        ANTENNAPARTIALMETALSIDEAREA 40.715  LAYER M3  ;
        ANTENNADIFFAREA 3.720  LAYER M2  ;
        ANTENNADIFFAREA 20.600  LAYER M3  ;
        ANTENNAPARTIALCUTAREA 0.135  LAYER V3  ;
        ANTENNAPARTIALCUTAREA 0.135  LAYER V2  ;
        PORT
        LAYER M2 ;
        RECT  36.370 249.580 37.100 250.000 ;
        LAYER M3 ;
        RECT  36.370 249.580 37.100 250.000 ;
        END
    END CIN
    PIN AVSSO
        DIRECTION INOUT ;
        USE ground ;
        PORT
        LAYER M2 ;
        RECT  0.000 147.040 65.000 154.520 ;
        LAYER M3 ;
        RECT  0.000 92.060 65.000 123.250 ;
        RECT  64.200 149.940 65.000 162.610 ;
        RECT  0.000 149.940 0.800 162.610 ;
        LAYER TOP_M ;
        RECT  0.000 92.060 65.000 123.250 ;
        RECT  0.000 155.410 65.000 162.610 ;
        END
    END AVSSO
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        PORT
        LAYER M3 ;
        RECT  64.200 130.680 65.000 140.840 ;
        RECT  0.000 130.680 0.800 140.840 ;
        LAYER TOP_M ;
        RECT  0.000 123.850 65.000 140.850 ;
        END
    END VSS
    PIN AVSS
        DIRECTION INOUT ;
        USE ground ;
        PORT
        LAYER M2 ;
        RECT  0.000 143.120 65.000 146.340 ;
        RECT  39.160 136.310 65.000 146.340 ;
        RECT  0.000 136.310 4.480 146.340 ;
        LAYER M3 ;
        RECT  64.200 141.450 65.000 148.880 ;
        RECT  0.000 141.450 0.800 148.880 ;
        LAYER TOP_M ;
        RECT  0.000 141.450 65.000 154.560 ;
        END
    END AVSS
    PIN AVDD
        DIRECTION INOUT ;
        USE power ;
        PORT
        LAYER M2 ;
        RECT  0.000 172.080 65.000 183.060 ;
        LAYER M3 ;
        RECT  64.200 163.510 65.000 190.890 ;
        RECT  0.000 163.510 0.800 190.890 ;
        LAYER TOP_M ;
        RECT  0.000 163.500 65.000 194.560 ;
        END
    END AVDD
    PIN AVDDO
        DIRECTION INOUT ;
        USE power ;
        PORT
        LAYER M2 ;
        RECT  0.000 186.470 65.000 194.870 ;
        LAYER M3 ;
        RECT  64.200 192.330 65.000 200.640 ;
        RECT  0.000 201.660 65.000 218.520 ;
        RECT  0.000 219.720 65.000 246.820 ;
        RECT  0.000 192.330 0.800 200.640 ;
        LAYER TOP_M ;
        RECT  0.000 195.170 65.000 200.640 ;
        RECT  0.000 201.660 65.000 221.520 ;
        RECT  0.000 222.720 65.000 246.820 ;
        END
    END AVDDO
    OBS
        LAYER M1 ;
        RECT  2.000 0.000 63.000 249.570 ;
        RECT  0.000 88.990 65.000 130.360 ;
        RECT  0.000 136.510 65.000 157.550 ;
        RECT  0.360 159.530 64.760 159.830 ;
        RECT  0.360 162.240 64.760 162.540 ;
        RECT  0.360 163.070 64.760 163.350 ;
        RECT  0.360 164.850 64.760 165.150 ;
        RECT  0.360 165.450 64.760 165.750 ;
        RECT  0.360 166.050 64.760 166.350 ;
        RECT  0.360 166.650 64.760 166.960 ;
        RECT  0.000 169.150 65.000 194.230 ;
        RECT  0.000 195.470 65.000 247.000 ;
        RECT  0.600 0.600 64.400 249.570 ;
        RECT  0.000 248.330 65.000 249.570 ;
        LAYER M2 ;
        RECT  12.700 195.440 14.380 249.400 ;
        RECT  50.010 195.470 52.040 249.400 ;
        RECT  0.600 195.660 64.400 241.930 ;
        RECT  35.160 195.660 64.400 248.790 ;
        RECT  0.600 195.660 31.560 249.400 ;
        RECT  35.160 195.660 35.580 249.400 ;
        RECT  37.890 195.660 64.400 249.400 ;
        RECT  3.940 195.660 7.950 249.570 ;
        RECT  18.470 183.720 52.450 185.680 ;
        RECT  0.600 183.850 64.400 185.680 ;
        RECT  44.225 183.850 54.190 185.870 ;
        RECT  55.120 183.850 63.815 185.870 ;
        RECT  52.275 155.260 52.595 171.290 ;
        RECT  53.375 155.210 54.975 171.290 ;
        RECT  0.600 155.310 64.400 171.290 ;
        RECT  26.590 155.310 26.910 171.455 ;
        RECT  24.140 155.310 25.740 171.470 ;
        RECT  23.040 155.310 23.360 171.475 ;
        RECT  58.240 155.310 58.520 171.480 ;
        RECT  2.000 0.000 63.000 60.210 ;
        RECT  0.600 0.600 64.400 60.210 ;
        RECT  0.600 0.600 1.210 135.520 ;
        RECT  0.600 91.020 64.400 135.520 ;
        RECT  4.070 91.020 60.930 135.690 ;
        RECT  5.270 91.020 38.370 142.330 ;
        RECT  5.415 136.510 38.560 142.520 ;
        LAYER M3 ;
        RECT  0.600 247.660 31.830 248.740 ;
        RECT  0.600 247.660 31.510 249.400 ;
        RECT  3.940 247.660 7.950 249.570 ;
        RECT  34.890 247.660 64.400 248.740 ;
        RECT  35.210 247.660 35.530 249.400 ;
        RECT  37.940 247.660 64.400 249.400 ;
        RECT  4.030 123.970 61.110 200.820 ;
        RECT  0.600 124.090 64.400 129.840 ;
        RECT  1.400 124.090 63.360 135.790 ;
        RECT  1.400 124.090 2.135 154.570 ;
        RECT  2.715 131.490 63.600 158.355 ;
        RECT  1.640 155.040 63.360 171.560 ;
        RECT  1.640 183.580 63.445 185.950 ;
        RECT  2.715 124.090 63.360 200.820 ;
        RECT  1.640 195.390 63.445 200.820 ;
        RECT  63.165 162.930 63.445 201.060 ;
        RECT  0.600 0.600 64.400 60.480 ;
        RECT  2.000 0.000 63.000 88.700 ;
        RECT  0.600 0.600 1.480 91.220 ;
        RECT  0.600 90.750 64.400 91.220 ;
        LAYER TOP_M ;
        RECT  0.600 247.690 64.400 248.850 ;
        RECT  0.600 247.690 31.620 249.400 ;
        RECT  35.100 247.690 35.640 249.400 ;
        RECT  37.830 247.690 64.400 249.400 ;
        RECT  2.000 0.000 63.000 91.190 ;
        RECT  0.600 0.600 64.400 91.190 ;
    END
END apc3d01

MACRO pfrelr
    CLASS ENDCAP BOTTOMRIGHT ;
    FOREIGN pfrelr 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 250.000 BY 250.000 ;
    SYMMETRY X Y R90 ;
    SITE CO_MSTR_c ;
    OBS
        LAYER M1 ;
        RECT  0.000 0.000 250.000 250.000 ;
        LAYER M2 ;
        RECT  0.000 0.000 250.000 250.000 ;
        LAYER M3 ;
        RECT  0.000 0.000 250.000 249.400 ;
        RECT  0.600 0.000 250.000 250.000 ;
        LAYER TOP_M ;
        RECT  0.000 0.000 250.000 249.400 ;
        RECT  0.600 0.000 250.000 250.000 ;
    END
END pfrelr

MACRO apfrelr
    CLASS ENDCAP BOTTOMRIGHT ;
    FOREIGN apfrelr 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 250.000 BY 250.000 ;
    SYMMETRY X Y R90 ;
    SITE CO_MSTR_c ;
    OBS
        LAYER M1 ;
        RECT  0.000 0.000 250.000 250.000 ;
        LAYER M2 ;
        RECT  0.000 0.000 250.000 250.000 ;
        LAYER M3 ;
        RECT  0.000 0.000 250.000 249.400 ;
        RECT  0.600 0.000 250.000 250.000 ;
        LAYER TOP_M ;
        RECT  0.000 0.000 250.000 249.400 ;
        RECT  0.600 0.000 250.000 250.000 ;
    END
END apfrelr

MACRO pfeedendringr
    CLASS PAD SPACER ;
    FOREIGN pfeedendringr 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.300 BY 250.000 ;
    SYMMETRY X Y R90 ;
    SITE IOSite_c ;
    OBS
        LAYER M1 ;
        RECT  0.000 0.000 1.300 250.000 ;
        LAYER M2 ;
        RECT  0.000 0.000 1.300 250.000 ;
        LAYER M3 ;
        RECT  0.000 0.000 1.300 250.000 ;
        LAYER TOP_M ;
        RECT  0.000 0.000 1.300 250.000 ;
    END
END pfeedendringr

MACRO pfeedendringl
    CLASS PAD SPACER ;
    FOREIGN pfeedendringl 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.300 BY 250.000 ;
    SYMMETRY X Y R90 ;
    SITE IOSite_c ;
    OBS
        LAYER M1 ;
        RECT  0.000 0.000 1.300 250.000 ;
        LAYER M2 ;
        RECT  0.000 0.000 1.300 250.000 ;
        LAYER M3 ;
        RECT  0.000 0.000 1.300 250.000 ;
        LAYER TOP_M ;
        RECT  0.000 0.000 1.300 250.000 ;
    END
END pfeedendringl

MACRO pfeed30000
    CLASS PAD SPACER ;
    FOREIGN pfeed30000 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 30.000 BY 250.000 ;
    SYMMETRY X Y R90 ;
    SITE IOSite_c ;
    OBS
        LAYER M1 ;
        RECT  0.000 0.000 30.000 250.000 ;
        LAYER M2 ;
        RECT  0.000 0.000 30.000 250.000 ;
        LAYER M3 ;
        RECT  0.000 0.000 30.000 250.000 ;
        LAYER TOP_M ;
        RECT  0.000 0.000 30.000 250.000 ;
    END
END pfeed30000

MACRO pfeed10000
    CLASS PAD SPACER ;
    FOREIGN pfeed10000 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.000 BY 250.000 ;
    SYMMETRY X Y R90 ;
    SITE IOSite_c ;
    OBS
        LAYER M1 ;
        RECT  0.000 0.000 10.000 250.000 ;
        LAYER M2 ;
        RECT  0.000 0.000 10.000 250.000 ;
        LAYER M3 ;
        RECT  0.000 0.000 10.000 250.000 ;
        LAYER TOP_M ;
        RECT  0.000 0.000 10.000 250.000 ;
    END
END pfeed10000

MACRO pfeed02000
    CLASS PAD SPACER ;
    FOREIGN pfeed02000 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.000 BY 250.000 ;
    SYMMETRY X Y R90 ;
    SITE IOSite_c ;
    OBS
        LAYER M1 ;
        RECT  0.000 0.000 2.000 250.000 ;
        LAYER M2 ;
        RECT  0.000 0.000 2.000 250.000 ;
        LAYER M3 ;
        RECT  0.000 0.000 2.000 250.000 ;
        LAYER TOP_M ;
        RECT  0.000 0.000 2.000 250.000 ;
    END
END pfeed02000

MACRO pfeed01000
    CLASS PAD SPACER ;
    FOREIGN pfeed01000 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.000 BY 250.000 ;
    SYMMETRY X Y R90 ;
    SITE IOSite_c ;
    OBS
        LAYER M1 ;
        RECT  0.000 0.000 1.000 250.000 ;
        LAYER M2 ;
        RECT  0.000 0.000 1.000 250.000 ;
        LAYER M3 ;
        RECT  0.000 0.000 1.000 250.000 ;
        LAYER TOP_M ;
        RECT  0.000 0.000 1.000 250.000 ;
    END
END pfeed01000

MACRO pfeed00540
    CLASS PAD SPACER ;
    FOREIGN pfeed00540 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.540 BY 250.000 ;
    SYMMETRY X Y R90 ;
    SITE IOSite_c ;
    OBS
        LAYER M1 ;
        RECT  0.000 0.000 0.540 250.000 ;
        LAYER M2 ;
        RECT  0.000 0.000 0.540 250.000 ;
        LAYER M3 ;
        RECT  0.000 0.000 0.540 250.000 ;
        LAYER TOP_M ;
        RECT  0.000 0.000 0.540 250.000 ;
    END
END pfeed00540

MACRO pfeed00120
    CLASS PAD SPACER ;
    FOREIGN pfeed00120 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.120 BY 250.000 ;
    SYMMETRY X Y R90 ;
    SITE IOSite_c ;
    OBS
        LAYER M1 ;
        RECT  0.000 0.000 0.120 250.000 ;
        LAYER M2 ;
        RECT  0.000 0.000 0.120 250.000 ;
        LAYER M3 ;
        RECT  0.000 0.000 0.120 250.000 ;
        LAYER TOP_M ;
        RECT  0.000 0.000 0.120 250.000 ;
    END
END pfeed00120

MACRO pfeed00040
    CLASS PAD SPACER ;
    FOREIGN pfeed00040 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.040 BY 250.000 ;
    SYMMETRY X Y R90 ;
    SITE IOSite_c ;
    OBS
        LAYER M1 ;
        RECT  0.000 0.000 0.040 250.000 ;
        LAYER M2 ;
        RECT  0.000 0.000 0.040 250.000 ;
        LAYER M3 ;
        RECT  0.000 0.000 0.040 250.000 ;
        LAYER TOP_M ;
        RECT  0.000 0.000 0.040 250.000 ;
    END
END pfeed00040

MACRO pfeed00010
    CLASS PAD SPACER ;
    FOREIGN pfeed00010 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.010 BY 250.000 ;
    SYMMETRY X Y R90 ;
    SITE IOSite_c ;
    OBS
        LAYER M1 ;
        RECT  0.000 0.000 0.010 250.000 ;
        LAYER M2 ;
        RECT  0.000 0.000 0.010 250.000 ;
        LAYER M3 ;
        RECT  0.000 0.000 0.010 250.000 ;
        LAYER TOP_M ;
        RECT  0.000 0.000 0.010 250.000 ;
    END
END pfeed00010

MACRO apfeedendringr
    CLASS PAD SPACER ;
    FOREIGN apfeedendringr 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 30.000 BY 250.000 ;
    SYMMETRY X Y R90 ;
    SITE IOSite_c ;
    OBS
        LAYER M1 ;
        RECT  0.000 0.000 30.000 250.000 ;
        LAYER M2 ;
        RECT  0.000 0.000 30.000 250.000 ;
        LAYER M3 ;
        RECT  0.000 0.000 30.000 250.000 ;
        LAYER TOP_M ;
        RECT  0.000 0.000 30.000 250.000 ;
    END
END apfeedendringr

MACRO apfeedendringl
    CLASS PAD SPACER ;
    FOREIGN apfeedendringl 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 30.000 BY 250.000 ;
    SYMMETRY X Y R90 ;
    SITE IOSite_c ;
    OBS
        LAYER M1 ;
        RECT  0.000 0.000 30.000 250.000 ;
        LAYER M2 ;
        RECT  0.000 0.000 30.000 250.000 ;
        LAYER M3 ;
        RECT  0.000 0.000 30.000 250.000 ;
        LAYER TOP_M ;
        RECT  0.000 0.000 30.000 250.000 ;
    END
END apfeedendringl

MACRO apfeed30000
    CLASS PAD SPACER ;
    FOREIGN apfeed30000 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 30.000 BY 250.000 ;
    SYMMETRY X Y R90 ;
    SITE IOSite_c ;
    OBS
        LAYER M1 ;
        RECT  0.000 0.000 30.000 250.000 ;
        LAYER M2 ;
        RECT  0.000 0.000 30.000 250.000 ;
        LAYER M3 ;
        RECT  0.000 0.000 30.000 250.000 ;
        LAYER TOP_M ;
        RECT  0.000 0.000 30.000 250.000 ;
    END
END apfeed30000

MACRO apfeed10000
    CLASS PAD SPACER ;
    FOREIGN apfeed10000 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.000 BY 250.000 ;
    SYMMETRY X Y R90 ;
    SITE IOSite_c ;
    OBS
        LAYER M1 ;
        RECT  0.000 0.000 10.000 250.000 ;
        LAYER M2 ;
        RECT  0.000 0.000 10.000 250.000 ;
        LAYER M3 ;
        RECT  0.000 0.000 10.000 250.000 ;
        LAYER TOP_M ;
        RECT  0.000 0.000 10.000 250.000 ;
    END
END apfeed10000

MACRO apfeed02000
    CLASS PAD SPACER ;
    FOREIGN apfeed02000 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.000 BY 250.000 ;
    SYMMETRY X Y R90 ;
    SITE IOSite_c ;
    OBS
        LAYER M1 ;
        RECT  0.000 0.000 2.000 250.000 ;
        LAYER M2 ;
        RECT  0.000 0.000 2.000 250.000 ;
        LAYER M3 ;
        RECT  0.000 0.000 2.000 250.000 ;
        LAYER TOP_M ;
        RECT  0.000 0.000 2.000 250.000 ;
    END
END apfeed02000

MACRO apfeed01000
    CLASS PAD SPACER ;
    FOREIGN apfeed01000 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.000 BY 250.000 ;
    SYMMETRY X Y R90 ;
    SITE IOSite_c ;
    OBS
        LAYER M1 ;
        RECT  0.000 0.000 1.000 250.000 ;
        LAYER M2 ;
        RECT  0.000 0.000 1.000 250.000 ;
        LAYER M3 ;
        RECT  0.000 0.000 1.000 250.000 ;
        LAYER TOP_M ;
        RECT  0.000 0.000 1.000 250.000 ;
    END
END apfeed01000

MACRO apfeed00540
    CLASS PAD SPACER ;
    FOREIGN apfeed00540 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.540 BY 250.000 ;
    SYMMETRY X Y R90 ;
    SITE IOSite_c ;
    OBS
        LAYER M1 ;
        RECT  0.000 0.000 0.540 250.000 ;
        LAYER M2 ;
        RECT  0.000 0.000 0.540 250.000 ;
        LAYER M3 ;
        RECT  0.000 0.000 0.540 250.000 ;
        LAYER TOP_M ;
        RECT  0.000 0.000 0.540 250.000 ;
    END
END apfeed00540

MACRO apfeed00120
    CLASS PAD SPACER ;
    FOREIGN apfeed00120 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.120 BY 250.000 ;
    SYMMETRY X Y R90 ;
    SITE IOSite_c ;
    OBS
        LAYER M1 ;
        RECT  0.000 0.000 0.120 250.000 ;
        LAYER M2 ;
        RECT  0.000 0.000 0.120 250.000 ;
        LAYER M3 ;
        RECT  0.000 0.000 0.120 250.000 ;
        LAYER TOP_M ;
        RECT  0.000 0.000 0.120 250.000 ;
    END
END apfeed00120

MACRO apfeed00040
    CLASS PAD SPACER ;
    FOREIGN apfeed00040 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.040 BY 250.000 ;
    SYMMETRY X Y R90 ;
    SITE IOSite_c ;
    OBS
        LAYER M1 ;
        RECT  0.000 0.000 0.040 250.000 ;
        LAYER M2 ;
        RECT  0.000 0.000 0.040 250.000 ;
        LAYER M3 ;
        RECT  0.000 0.000 0.040 250.000 ;
        LAYER TOP_M ;
        RECT  0.000 0.000 0.040 250.000 ;
    END
END apfeed00040

MACRO apfeed00010
    CLASS PAD SPACER ;
    FOREIGN apfeed00010 0 0 ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.010 BY 250.000 ;
    SYMMETRY X Y R90 ;
    SITE IOSite_c ;
    OBS
        LAYER M1 ;
        RECT  0.000 0.000 0.010 250.000 ;
        LAYER M2 ;
        RECT  0.000 0.000 0.010 250.000 ;
        LAYER M3 ;
        RECT  0.000 0.000 0.010 250.000 ;
        LAYER TOP_M ;
        RECT  0.000 0.000 0.010 250.000 ;
    END
END apfeed00010

END LIBRARY
